
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_register_file_WORD_SIZE32_ADDR_SIZE5 is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_register_file_WORD_SIZE32_ADDR_SIZE5;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_register_file_WORD_SIZE32_ADDR_SIZE5.all;

entity register_file_WORD_SIZE32_ADDR_SIZE5 is

   port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
         ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
         std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector (31
         downto 0));

end register_file_WORD_SIZE32_ADDR_SIZE5;

architecture SYN_Beh of register_file_WORD_SIZE32_ADDR_SIZE5 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
      n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, 
      n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, 
      n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, 
      n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, 
      n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, 
      n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, 
      n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, 
      n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, 
      n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, 
      n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, 
      n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, 
      n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, 
      n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, 
      n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, 
      n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, 
      n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, 
      n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, 
      n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, 
      n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, 
      n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, 
      n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, 
      n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, 
      n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, 
      n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, 
      n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, 
      n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, 
      n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, 
      n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, 
      n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, 
      n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, 
      n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, 
      n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, 
      n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, 
      n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, 
      n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, 
      n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, 
      n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, 
      n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, 
      n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, 
      n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, 
      n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, 
      n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, 
      n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, 
      n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, 
      n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, 
      n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, 
      n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, 
      n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, 
      n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, 
      n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, 
      n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, 
      n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, 
      n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, 
      n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, 
      n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, 
      n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, 
      n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, 
      n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, 
      n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, 
      n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, 
      n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, 
      n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, 
      n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, 
      n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, 
      n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, 
      n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, 
      n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, 
      n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, 
      n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, 
      n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, 
      n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, 
      n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, 
      n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, 
      n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, 
      n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, 
      n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, 
      n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, 
      n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, 
      n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, 
      n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, 
      n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, 
      n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, 
      n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, 
      n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, 
      n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, 
      n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, 
      n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, 
      n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, 
      n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, 
      n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, 
      n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, 
      n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, 
      n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, 
      n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, 
      n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, 
      n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, 
      n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, 
      n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, 
      n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, 
      n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, 
      n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, 
      n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, 
      n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, 
      n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, 
      n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, 
      n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, 
      n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, 
      n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n8988, n8989, 
      n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, 
      n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, 
      n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, 
      n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, 
      n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, 
      n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, 
      n9146, n9147, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, 
      n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, 
      n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, 
      n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, 
      n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, 
      n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, 
      n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, 
      n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, 
      n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, 
      n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, 
      n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, 
      n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, 
      n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, 
      n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, 
      n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, 
      n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, 
      n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, 
      n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, 
      n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, 
      n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, 
      n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, 
      n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, 
      n9622, n9623, n9624, n9625, n9626, n9627, n9630, n9631, n9632, n9633, 
      n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, 
      n9644, n9645, n9646, n9647, n9648, n9659, n9670, n9671, n9672, n9673, 
      n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, 
      n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, 
      n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9893, n9895, 
      n9897, n9899, n9901, n9903, n9905, n9907, n9909, n9911, n9913, n9915, 
      n9917, n9919, n9921, n9923, n9925, n9927, n9929, n9931, n9933, n9935, 
      n9937, n9939, n9941, n9943, n9945, n9947, n9949, n9951, n9953, n9955, 
      n10986, n10987, n10988, n10989, n10990, n10991, n10996, n10997, n10998, 
      n10999, n11004, n11005, n11006, n11007, n11948, n11949, n11950, n11951, 
      n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960, 
      n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969, 
      n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978, 
      n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987, 
      n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995, n11996, 
      n11997, n11998, n11999, n12000, n12001, n12002, n12003, n12004, n12005, 
      n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013, n12014, 
      n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023, 
      n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032, 
      n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12042, n12043, 
      n12044, n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054, 
      n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063, 
      n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072, 
      n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081, 
      n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090, 
      n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099, 
      n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107, n12108, 
      n12109, n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117, 
      n12118, n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126, 
      n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135, 
      n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144, 
      n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153, 
      n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162, 
      n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171, 
      n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179, n12180, 
      n12181, n12182, n12183, n12184, n12185, n12186, n12187, n12188, n12189, 
      n12190, n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198, 
      n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207, 
      n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216, 
      n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225, 
      n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234, 
      n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243, 
      n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251, n12252, 
      n12253, n12254, n12255, n12256, n12257, n12258, n12259, n12260, n12261, 
      n12262, n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270, 
      n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279, 
      n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288, 
      n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297, 
      n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306, 
      n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315, 
      n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323, n12324, 
      n12325, n12326, n12327, n12328, n12329, n12330, n12331, n12332, n12333, 
      n12334, n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342, 
      n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351, 
      n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360, 
      n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369, 
      n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378, 
      n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387, 
      n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396, 
      n12397, n12398, n12399, n12400, n12401, n12402, n12403, n12404, n12405, 
      n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414, 
      n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423, 
      n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432, 
      n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441, 
      n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450, 
      n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459, 
      n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468, 
      n12469, n12470, n12471, n12472, n12473, n12474, n12475, n12476, n12477, 
      n12478, n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486, 
      n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495, 
      n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504, 
      n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513, 
      n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522, 
      n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531, 
      n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539, n12540, 
      n12541, n12542, n12543, n12544, n12545, n12546, n12547, n12548, n12549, 
      n12550, n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558, 
      n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567, 
      n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576, 
      n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585, 
      n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594, 
      n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603, 
      n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611, n12612, 
      n12613, n12614, n12615, n12616, n12617, n12618, n12619, n12620, n12623, 
      n12624, n12625, n12628, n12629, n12630, n12631, n12632, n12633, n12634, 
      n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643, 
      n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652, 
      n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12660, n12661, 
      n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670, 
      n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679, 
      n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688, 
      n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697, 
      n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706, 
      n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715, 
      n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724, 
      n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732, n12733, 
      n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742, 
      n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751, 
      n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760, 
      n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769, 
      n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778, 
      n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787, 
      n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796, 
      n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805, 
      n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814, 
      n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823, 
      n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832, 
      n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841, 
      n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850, 
      n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859, 
      n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868, 
      n12869, n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877, 
      n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886, 
      n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895, 
      n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904, 
      n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913, 
      n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922, 
      n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931, 
      n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940, 
      n12941, n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949, 
      n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958, 
      n12959, n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967, 
      n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976, 
      n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985, 
      n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994, 
      n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003, 
      n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011, n13012, 
      n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021, 
      n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030, 
      n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039, 
      n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048, 
      n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057, 
      n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066, 
      n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075, 
      n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084, 
      n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093, 
      n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102, 
      n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111, 
      n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120, 
      n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129, 
      n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138, 
      n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147, 
      n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156, 
      n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165, 
      n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174, 
      n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183, 
      n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192, 
      n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201, 
      n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210, 
      n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219, 
      n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228, 
      n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237, 
      n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246, 
      n13247, n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255, 
      n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264, 
      n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273, 
      n13274, n13275, n13300, n13301, n13302, n13303, n13304, n13305, n13306, 
      n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315, 
      n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13348, 
      n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357, 
      n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366, 
      n13367, n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375, 
      n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384, 
      n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393, 
      n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402, 
      n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411, 
      n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419, n13492, 
      n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501, 
      n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509, n13510, 
      n13511, n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519, 
      n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528, 
      n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537, 
      n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546, 
      n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555, 
      n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13636, 
      n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645, 
      n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653, n13654, 
      n13655, n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663, 
      n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672, 
      n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681, 
      n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690, 
      n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699, 
      n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707, n13708, 
      n13709, n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717, 
      n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725, n13726, 
      n13727, n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735, 
      n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744, 
      n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753, 
      n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762, 
      n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771, 
      n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779, n13780, 
      n13781, n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789, 
      n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797, n13798, 
      n13799, n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807, 
      n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816, 
      n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825, 
      n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834, 
      n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843, 
      n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851, n13852, 
      n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861, 
      n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869, n13870, 
      n13871, n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879, 
      n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888, 
      n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897, 
      n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906, 
      n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915, 
      n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923, n13924, 
      n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933, 
      n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941, n13942, 
      n13943, n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951, 
      n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960, 
      n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969, 
      n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978, 
      n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987, 
      n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995, n13996, 
      n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005, 
      n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013, n14014, 
      n14015, n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023, 
      n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032, 
      n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041, 
      n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050, 
      n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059, 
      n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068, 
      n14069, n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077, 
      n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085, n14086, 
      n14087, n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095, 
      n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104, 
      n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113, 
      n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122, 
      n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131, 
      n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140, 
      n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149, 
      n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157, n14158, 
      n14159, n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167, 
      n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176, 
      n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185, 
      n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194, 
      n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203, 
      n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211, n14212, 
      n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221, 
      n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229, n14230, 
      n14231, n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239, 
      n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248, 
      n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257, 
      n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266, 
      n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275, 
      n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284, 
      n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293, 
      n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301, n14302, 
      n14303, n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311, 
      n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320, 
      n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329, 
      n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338, 
      n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347, 
      n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355, n14356, 
      n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365, 
      n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373, n14374, 
      n14375, n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383, 
      n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392, 
      n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401, 
      n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410, 
      n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419, 
      n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428, 
      n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437, 
      n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445, n14446, 
      n14447, n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455, 
      n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464, 
      n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473, 
      n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482, 
      n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491, 
      n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500, 
      n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509, 
      n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517, n14518, 
      n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527, 
      n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536, 
      n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545, 
      n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554, 
      n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563, 
      n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571, n14572, 
      n14573, n14574, n14575, n14576, n14577, n14578, n14579, n14580, n14581, 
      n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589, n14590, 
      n14591, n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599, 
      n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608, 
      n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617, 
      n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626, 
      n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635, 
      n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644, 
      n14645, n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653, 
      n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661, n14662, 
      n14663, n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671, 
      n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680, 
      n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689, 
      n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698, 
      n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707, 
      n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715, n14716, 
      n14717, n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725, 
      n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14733, n14734, 
      n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743, 
      n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752, 
      n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761, 
      n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770, 
      n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779, 
      n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787, n14788, 
      n14789, n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797, 
      n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805, n14806, 
      n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815, 
      n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824, 
      n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833, 
      n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842, 
      n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851, 
      n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859, n14860, 
      n14861, n14862, n14863, n14864, n14865, n14866, n14867, n14868, n14869, 
      n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877, n14878, 
      n14879, n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887, 
      n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896, 
      n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905, 
      n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914, 
      n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923, 
      n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931, n14932, 
      n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940, n14941, 
      n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949, n14950, 
      n14951, n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14959, 
      n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968, 
      n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977, 
      n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986, 
      n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995, 
      n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003, n15004, 
      n15005, n15006, n15007, n15008, n15009, n15010, n15011, n15012, n15013, 
      n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021, n15022, 
      n15023, n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031, 
      n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040, 
      n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049, 
      n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058, 
      n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067, 
      n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075, n15076, 
      n15077, n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085, 
      n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093, n15094, 
      n15095, n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103, 
      n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112, 
      n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121, 
      n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130, 
      n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139, 
      n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147, n15148, 
      n15149, n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157, 
      n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165, n15166, 
      n15167, n15168, n15169, n15170, n15171, n_1000, n_1001, n_1002, n_1003, 
      n_1004, n_1005, n_1006, n_1007, n_1008, n_1009, n_1010, n_1011, n_1012, 
      n_1013, n_1014, n_1015, n_1016, n_1017, n_1018, n_1019, n_1020, n_1021, 
      n_1022, n_1023, n_1024, n_1025, n_1026, n_1027, n_1028, n_1029, n_1030, 
      n_1031, n_1032, n_1033, n_1034, n_1035, n_1036, n_1037, n_1038, n_1039, 
      n_1040, n_1041, n_1042, n_1043, n_1044, n_1045, n_1046, n_1047, n_1048, 
      n_1049, n_1050, n_1051, n_1052, n_1053, n_1054, n_1055, n_1056, n_1057, 
      n_1058, n_1059, n_1060, n_1061, n_1062, n_1063, n_1064, n_1065, n_1066, 
      n_1067, n_1068, n_1069, n_1070, n_1071, n_1072, n_1073, n_1074, n_1075, 
      n_1076, n_1077, n_1078, n_1079, n_1080, n_1081, n_1082, n_1083, n_1084, 
      n_1085, n_1086, n_1087, n_1088, n_1089, n_1090, n_1091, n_1092, n_1093, 
      n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, n_1100, n_1101, n_1102, 
      n_1103, n_1104, n_1105, n_1106, n_1107, n_1108, n_1109, n_1110, n_1111, 
      n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, n_1119, n_1120, 
      n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, n_1127, n_1128, n_1129, 
      n_1130, n_1131, n_1132, n_1133, n_1134, n_1135, n_1136, n_1137, n_1138, 
      n_1139, n_1140, n_1141, n_1142, n_1143, n_1144, n_1145, n_1146, n_1147, 
      n_1148, n_1149, n_1150, n_1151, n_1152, n_1153, n_1154, n_1155, n_1156, 
      n_1157, n_1158, n_1159, n_1160, n_1161, n_1162, n_1163, n_1164, n_1165, 
      n_1166, n_1167, n_1168, n_1169, n_1170, n_1171, n_1172, n_1173, n_1174, 
      n_1175, n_1176, n_1177, n_1178, n_1179, n_1180, n_1181, n_1182, n_1183, 
      n_1184, n_1185, n_1186, n_1187, n_1188, n_1189, n_1190, n_1191, n_1192, 
      n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, n_1199, n_1200, n_1201, 
      n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, n_1208, n_1209, n_1210, 
      n_1211, n_1212, n_1213, n_1214, n_1215, n_1216, n_1217, n_1218, n_1219, 
      n_1220, n_1221, n_1222, n_1223, n_1224, n_1225, n_1226, n_1227, n_1228, 
      n_1229, n_1230, n_1231, n_1232, n_1233, n_1234, n_1235, n_1236, n_1237, 
      n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, n_1244, n_1245, n_1246, 
      n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, n_1253, n_1254, n_1255, 
      n_1256, n_1257, n_1258, n_1259, n_1260, n_1261, n_1262, n_1263, n_1264, 
      n_1265, n_1266, n_1267, n_1268, n_1269, n_1270, n_1271, n_1272, n_1273, 
      n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, n_1280, n_1281, n_1282, 
      n_1283, n_1284, n_1285, n_1286, n_1287, n_1288, n_1289, n_1290, n_1291, 
      n_1292, n_1293, n_1294, n_1295, n_1296, n_1297, n_1298, n_1299, n_1300, 
      n_1301, n_1302, n_1303, n_1304, n_1305, n_1306, n_1307, n_1308, n_1309, 
      n_1310, n_1311, n_1312, n_1313, n_1314, n_1315, n_1316, n_1317, n_1318, 
      n_1319, n_1320, n_1321, n_1322, n_1323, n_1324, n_1325, n_1326, n_1327, 
      n_1328, n_1329, n_1330, n_1331, n_1332, n_1333, n_1334, n_1335, n_1336, 
      n_1337, n_1338, n_1339, n_1340, n_1341, n_1342, n_1343, n_1344, n_1345, 
      n_1346, n_1347, n_1348, n_1349, n_1350, n_1351, n_1352, n_1353, n_1354, 
      n_1355, n_1356, n_1357, n_1358, n_1359, n_1360, n_1361, n_1362, n_1363, 
      n_1364, n_1365, n_1366, n_1367, n_1368, n_1369, n_1370, n_1371, n_1372, 
      n_1373, n_1374, n_1375, n_1376, n_1377, n_1378, n_1379, n_1380, n_1381, 
      n_1382, n_1383, n_1384, n_1385, n_1386, n_1387, n_1388, n_1389, n_1390, 
      n_1391, n_1392, n_1393, n_1394, n_1395, n_1396, n_1397, n_1398, n_1399, 
      n_1400, n_1401, n_1402, n_1403, n_1404, n_1405, n_1406, n_1407, n_1408, 
      n_1409, n_1410, n_1411, n_1412, n_1413, n_1414, n_1415, n_1416, n_1417, 
      n_1418, n_1419, n_1420, n_1421, n_1422, n_1423, n_1424, n_1425, n_1426, 
      n_1427, n_1428, n_1429, n_1430, n_1431, n_1432, n_1433, n_1434, n_1435, 
      n_1436, n_1437, n_1438, n_1439, n_1440, n_1441, n_1442, n_1443, n_1444, 
      n_1445, n_1446, n_1447, n_1448, n_1449, n_1450, n_1451, n_1452, n_1453, 
      n_1454, n_1455, n_1456, n_1457, n_1458, n_1459, n_1460, n_1461, n_1462, 
      n_1463, n_1464, n_1465, n_1466, n_1467, n_1468, n_1469, n_1470, n_1471, 
      n_1472, n_1473, n_1474, n_1475, n_1476, n_1477, n_1478, n_1479, n_1480, 
      n_1481, n_1482, n_1483, n_1484, n_1485, n_1486, n_1487, n_1488, n_1489, 
      n_1490, n_1491, n_1492, n_1493, n_1494, n_1495, n_1496, n_1497, n_1498, 
      n_1499, n_1500, n_1501, n_1502, n_1503, n_1504, n_1505, n_1506, n_1507, 
      n_1508, n_1509, n_1510, n_1511, n_1512, n_1513, n_1514, n_1515, n_1516, 
      n_1517, n_1518, n_1519, n_1520, n_1521, n_1522, n_1523, n_1524, n_1525, 
      n_1526, n_1527, n_1528, n_1529, n_1530, n_1531, n_1532, n_1533, n_1534, 
      n_1535, n_1536, n_1537, n_1538, n_1539, n_1540, n_1541, n_1542, n_1543 : 
      std_logic;

begin
   
   REGISTERS_reg_0_31_inst : DFF_X1 port map( D => n2365, CK => CLK, Q => 
                           n_1000, QN => n13767);
   REGISTERS_reg_0_30_inst : DFF_X1 port map( D => n2364, CK => CLK, Q => 
                           n_1001, QN => n13766);
   REGISTERS_reg_0_29_inst : DFF_X1 port map( D => n2363, CK => CLK, Q => 
                           n_1002, QN => n13765);
   REGISTERS_reg_0_28_inst : DFF_X1 port map( D => n2362, CK => CLK, Q => 
                           n_1003, QN => n13764);
   REGISTERS_reg_0_27_inst : DFF_X1 port map( D => n2361, CK => CLK, Q => 
                           n_1004, QN => n13763);
   REGISTERS_reg_0_26_inst : DFF_X1 port map( D => n2360, CK => CLK, Q => 
                           n_1005, QN => n13762);
   REGISTERS_reg_0_25_inst : DFF_X1 port map( D => n2359, CK => CLK, Q => 
                           n_1006, QN => n13761);
   REGISTERS_reg_0_24_inst : DFF_X1 port map( D => n2358, CK => CLK, Q => 
                           n_1007, QN => n13760);
   REGISTERS_reg_0_23_inst : DFF_X1 port map( D => n2357, CK => CLK, Q => 
                           n_1008, QN => n13791);
   REGISTERS_reg_0_22_inst : DFF_X1 port map( D => n2356, CK => CLK, Q => 
                           n_1009, QN => n13790);
   REGISTERS_reg_0_21_inst : DFF_X1 port map( D => n2355, CK => CLK, Q => 
                           n_1010, QN => n13789);
   REGISTERS_reg_0_20_inst : DFF_X1 port map( D => n2354, CK => CLK, Q => 
                           n_1011, QN => n13788);
   REGISTERS_reg_0_19_inst : DFF_X1 port map( D => n2353, CK => CLK, Q => 
                           n_1012, QN => n13787);
   REGISTERS_reg_0_18_inst : DFF_X1 port map( D => n2352, CK => CLK, Q => 
                           n_1013, QN => n13786);
   REGISTERS_reg_0_17_inst : DFF_X1 port map( D => n2351, CK => CLK, Q => 
                           n_1014, QN => n13785);
   REGISTERS_reg_0_16_inst : DFF_X1 port map( D => n2350, CK => CLK, Q => 
                           n_1015, QN => n13784);
   REGISTERS_reg_0_15_inst : DFF_X1 port map( D => n2349, CK => CLK, Q => 
                           n_1016, QN => n13783);
   REGISTERS_reg_0_14_inst : DFF_X1 port map( D => n2348, CK => CLK, Q => 
                           n_1017, QN => n13782);
   REGISTERS_reg_0_13_inst : DFF_X1 port map( D => n2347, CK => CLK, Q => 
                           n_1018, QN => n13781);
   REGISTERS_reg_0_12_inst : DFF_X1 port map( D => n2346, CK => CLK, Q => 
                           n_1019, QN => n13780);
   REGISTERS_reg_0_11_inst : DFF_X1 port map( D => n2345, CK => CLK, Q => 
                           n_1020, QN => n13855);
   REGISTERS_reg_0_10_inst : DFF_X1 port map( D => n2344, CK => CLK, Q => 
                           n_1021, QN => n13854);
   REGISTERS_reg_0_9_inst : DFF_X1 port map( D => n2343, CK => CLK, Q => n_1022
                           , QN => n13853);
   REGISTERS_reg_0_8_inst : DFF_X1 port map( D => n2342, CK => CLK, Q => n_1023
                           , QN => n13852);
   REGISTERS_reg_0_7_inst : DFF_X1 port map( D => n2341, CK => CLK, Q => n_1024
                           , QN => n13851);
   REGISTERS_reg_0_6_inst : DFF_X1 port map( D => n2340, CK => CLK, Q => n_1025
                           , QN => n13850);
   REGISTERS_reg_0_5_inst : DFF_X1 port map( D => n2339, CK => CLK, Q => n_1026
                           , QN => n13849);
   REGISTERS_reg_0_4_inst : DFF_X1 port map( D => n2338, CK => CLK, Q => n_1027
                           , QN => n13848);
   REGISTERS_reg_0_3_inst : DFF_X1 port map( D => n2337, CK => CLK, Q => n_1028
                           , QN => n13847);
   REGISTERS_reg_0_2_inst : DFF_X1 port map( D => n2336, CK => CLK, Q => n_1029
                           , QN => n13846);
   REGISTERS_reg_0_1_inst : DFF_X1 port map( D => n2335, CK => CLK, Q => n_1030
                           , QN => n13845);
   REGISTERS_reg_0_0_inst : DFF_X1 port map( D => n2334, CK => CLK, Q => n_1031
                           , QN => n13844);
   REGISTERS_reg_1_31_inst : DFF_X1 port map( D => n2333, CK => CLK, Q => 
                           n_1032, QN => n13871);
   REGISTERS_reg_1_30_inst : DFF_X1 port map( D => n2332, CK => CLK, Q => 
                           n_1033, QN => n13870);
   REGISTERS_reg_1_29_inst : DFF_X1 port map( D => n2331, CK => CLK, Q => 
                           n_1034, QN => n13869);
   REGISTERS_reg_1_28_inst : DFF_X1 port map( D => n2330, CK => CLK, Q => 
                           n_1035, QN => n13868);
   REGISTERS_reg_1_27_inst : DFF_X1 port map( D => n2329, CK => CLK, Q => 
                           n_1036, QN => n13867);
   REGISTERS_reg_1_26_inst : DFF_X1 port map( D => n2328, CK => CLK, Q => 
                           n_1037, QN => n13866);
   REGISTERS_reg_1_25_inst : DFF_X1 port map( D => n2327, CK => CLK, Q => 
                           n_1038, QN => n13865);
   REGISTERS_reg_1_24_inst : DFF_X1 port map( D => n2326, CK => CLK, Q => 
                           n_1039, QN => n13864);
   REGISTERS_reg_1_23_inst : DFF_X1 port map( D => n2325, CK => CLK, Q => 
                           n_1040, QN => n14141);
   REGISTERS_reg_1_22_inst : DFF_X1 port map( D => n2324, CK => CLK, Q => 
                           n_1041, QN => n14140);
   REGISTERS_reg_1_21_inst : DFF_X1 port map( D => n2323, CK => CLK, Q => 
                           n_1042, QN => n14139);
   REGISTERS_reg_1_20_inst : DFF_X1 port map( D => n2322, CK => CLK, Q => 
                           n_1043, QN => n14138);
   REGISTERS_reg_1_19_inst : DFF_X1 port map( D => n2321, CK => CLK, Q => 
                           n_1044, QN => n14137);
   REGISTERS_reg_1_18_inst : DFF_X1 port map( D => n2320, CK => CLK, Q => 
                           n_1045, QN => n14136);
   REGISTERS_reg_1_17_inst : DFF_X1 port map( D => n2319, CK => CLK, Q => 
                           n_1046, QN => n14135);
   REGISTERS_reg_1_16_inst : DFF_X1 port map( D => n2318, CK => CLK, Q => 
                           n_1047, QN => n14134);
   REGISTERS_reg_1_15_inst : DFF_X1 port map( D => n2317, CK => CLK, Q => 
                           n_1048, QN => n14133);
   REGISTERS_reg_1_14_inst : DFF_X1 port map( D => n2316, CK => CLK, Q => 
                           n_1049, QN => n14132);
   REGISTERS_reg_1_13_inst : DFF_X1 port map( D => n2315, CK => CLK, Q => 
                           n_1050, QN => n14131);
   REGISTERS_reg_1_12_inst : DFF_X1 port map( D => n2314, CK => CLK, Q => 
                           n_1051, QN => n14130);
   REGISTERS_reg_1_11_inst : DFF_X1 port map( D => n2313, CK => CLK, Q => 
                           n_1052, QN => n14129);
   REGISTERS_reg_1_10_inst : DFF_X1 port map( D => n2312, CK => CLK, Q => 
                           n_1053, QN => n14128);
   REGISTERS_reg_1_9_inst : DFF_X1 port map( D => n2311, CK => CLK, Q => n_1054
                           , QN => n14127);
   REGISTERS_reg_1_8_inst : DFF_X1 port map( D => n2310, CK => CLK, Q => n_1055
                           , QN => n14126);
   REGISTERS_reg_1_7_inst : DFF_X1 port map( D => n2309, CK => CLK, Q => n_1056
                           , QN => n14125);
   REGISTERS_reg_1_6_inst : DFF_X1 port map( D => n2308, CK => CLK, Q => n_1057
                           , QN => n14124);
   REGISTERS_reg_1_5_inst : DFF_X1 port map( D => n2307, CK => CLK, Q => n_1058
                           , QN => n14123);
   REGISTERS_reg_1_4_inst : DFF_X1 port map( D => n2306, CK => CLK, Q => n_1059
                           , QN => n14122);
   REGISTERS_reg_1_3_inst : DFF_X1 port map( D => n2305, CK => CLK, Q => n_1060
                           , QN => n14121);
   REGISTERS_reg_1_2_inst : DFF_X1 port map( D => n2304, CK => CLK, Q => n_1061
                           , QN => n14120);
   REGISTERS_reg_1_1_inst : DFF_X1 port map( D => n2303, CK => CLK, Q => n_1062
                           , QN => n14119);
   REGISTERS_reg_1_0_inst : DFF_X1 port map( D => n2302, CK => CLK, Q => n_1063
                           , QN => n14118);
   REGISTERS_reg_2_31_inst : DFF_X1 port map( D => n2301, CK => CLK, Q => 
                           n_1064, QN => n13831);
   REGISTERS_reg_2_30_inst : DFF_X1 port map( D => n2300, CK => CLK, Q => 
                           n_1065, QN => n13830);
   REGISTERS_reg_2_29_inst : DFF_X1 port map( D => n2299, CK => CLK, Q => 
                           n_1066, QN => n13829);
   REGISTERS_reg_2_28_inst : DFF_X1 port map( D => n2298, CK => CLK, Q => 
                           n_1067, QN => n13828);
   REGISTERS_reg_2_27_inst : DFF_X1 port map( D => n2297, CK => CLK, Q => 
                           n_1068, QN => n13827);
   REGISTERS_reg_2_26_inst : DFF_X1 port map( D => n2296, CK => CLK, Q => 
                           n_1069, QN => n13826);
   REGISTERS_reg_2_25_inst : DFF_X1 port map( D => n2295, CK => CLK, Q => 
                           n_1070, QN => n13825);
   REGISTERS_reg_2_24_inst : DFF_X1 port map( D => n2294, CK => CLK, Q => 
                           n_1071, QN => n13824);
   REGISTERS_reg_2_23_inst : DFF_X1 port map( D => n2293, CK => CLK, Q => 
                           n_1072, QN => n14085);
   REGISTERS_reg_2_22_inst : DFF_X1 port map( D => n2292, CK => CLK, Q => 
                           n_1073, QN => n14084);
   REGISTERS_reg_2_21_inst : DFF_X1 port map( D => n2291, CK => CLK, Q => 
                           n_1074, QN => n14083);
   REGISTERS_reg_2_20_inst : DFF_X1 port map( D => n2290, CK => CLK, Q => 
                           n_1075, QN => n14082);
   REGISTERS_reg_2_19_inst : DFF_X1 port map( D => n2289, CK => CLK, Q => 
                           n_1076, QN => n14081);
   REGISTERS_reg_2_18_inst : DFF_X1 port map( D => n2288, CK => CLK, Q => 
                           n_1077, QN => n14080);
   REGISTERS_reg_2_17_inst : DFF_X1 port map( D => n2287, CK => CLK, Q => 
                           n_1078, QN => n14079);
   REGISTERS_reg_2_16_inst : DFF_X1 port map( D => n2286, CK => CLK, Q => 
                           n_1079, QN => n14078);
   REGISTERS_reg_2_15_inst : DFF_X1 port map( D => n2285, CK => CLK, Q => 
                           n_1080, QN => n14077);
   REGISTERS_reg_2_14_inst : DFF_X1 port map( D => n2284, CK => CLK, Q => 
                           n_1081, QN => n14076);
   REGISTERS_reg_2_13_inst : DFF_X1 port map( D => n2283, CK => CLK, Q => 
                           n_1082, QN => n14075);
   REGISTERS_reg_2_12_inst : DFF_X1 port map( D => n2282, CK => CLK, Q => 
                           n_1083, QN => n14074);
   REGISTERS_reg_2_11_inst : DFF_X1 port map( D => n2281, CK => CLK, Q => 
                           n_1084, QN => n14073);
   REGISTERS_reg_2_10_inst : DFF_X1 port map( D => n2280, CK => CLK, Q => 
                           n_1085, QN => n14072);
   REGISTERS_reg_2_9_inst : DFF_X1 port map( D => n2279, CK => CLK, Q => n_1086
                           , QN => n14071);
   REGISTERS_reg_2_8_inst : DFF_X1 port map( D => n2278, CK => CLK, Q => n_1087
                           , QN => n14070);
   REGISTERS_reg_2_7_inst : DFF_X1 port map( D => n2277, CK => CLK, Q => n_1088
                           , QN => n14093);
   REGISTERS_reg_2_6_inst : DFF_X1 port map( D => n2276, CK => CLK, Q => n_1089
                           , QN => n14092);
   REGISTERS_reg_2_5_inst : DFF_X1 port map( D => n2275, CK => CLK, Q => n_1090
                           , QN => n14091);
   REGISTERS_reg_2_4_inst : DFF_X1 port map( D => n2274, CK => CLK, Q => n_1091
                           , QN => n14090);
   REGISTERS_reg_2_3_inst : DFF_X1 port map( D => n2273, CK => CLK, Q => n_1092
                           , QN => n14089);
   REGISTERS_reg_2_2_inst : DFF_X1 port map( D => n2272, CK => CLK, Q => n_1093
                           , QN => n14088);
   REGISTERS_reg_2_1_inst : DFF_X1 port map( D => n2271, CK => CLK, Q => n_1094
                           , QN => n14087);
   REGISTERS_reg_2_0_inst : DFF_X1 port map( D => n2270, CK => CLK, Q => n_1095
                           , QN => n14086);
   REGISTERS_reg_3_31_inst : DFF_X1 port map( D => n2269, CK => CLK, Q => n9701
                           , QN => n14011);
   REGISTERS_reg_3_30_inst : DFF_X1 port map( D => n2268, CK => CLK, Q => n9700
                           , QN => n14010);
   REGISTERS_reg_3_29_inst : DFF_X1 port map( D => n2267, CK => CLK, Q => n9699
                           , QN => n14009);
   REGISTERS_reg_3_28_inst : DFF_X1 port map( D => n2266, CK => CLK, Q => n9698
                           , QN => n14008);
   REGISTERS_reg_3_27_inst : DFF_X1 port map( D => n2265, CK => CLK, Q => n9697
                           , QN => n14007);
   REGISTERS_reg_3_26_inst : DFF_X1 port map( D => n2264, CK => CLK, Q => n9696
                           , QN => n14006);
   REGISTERS_reg_3_25_inst : DFF_X1 port map( D => n2263, CK => CLK, Q => n9695
                           , QN => n14005);
   REGISTERS_reg_3_24_inst : DFF_X1 port map( D => n2262, CK => CLK, Q => n9694
                           , QN => n14004);
   REGISTERS_reg_3_23_inst : DFF_X1 port map( D => n2261, CK => CLK, Q => n9693
                           , QN => n14481);
   REGISTERS_reg_3_22_inst : DFF_X1 port map( D => n2260, CK => CLK, Q => n9692
                           , QN => n14480);
   REGISTERS_reg_3_21_inst : DFF_X1 port map( D => n2259, CK => CLK, Q => n9691
                           , QN => n14479);
   REGISTERS_reg_3_20_inst : DFF_X1 port map( D => n2258, CK => CLK, Q => n9690
                           , QN => n14478);
   REGISTERS_reg_3_19_inst : DFF_X1 port map( D => n2257, CK => CLK, Q => n9689
                           , QN => n14477);
   REGISTERS_reg_3_18_inst : DFF_X1 port map( D => n2256, CK => CLK, Q => n9688
                           , QN => n14476);
   REGISTERS_reg_3_17_inst : DFF_X1 port map( D => n2255, CK => CLK, Q => n9687
                           , QN => n14475);
   REGISTERS_reg_3_16_inst : DFF_X1 port map( D => n2254, CK => CLK, Q => n9686
                           , QN => n14474);
   REGISTERS_reg_3_15_inst : DFF_X1 port map( D => n2253, CK => CLK, Q => n9685
                           , QN => n14473);
   REGISTERS_reg_3_14_inst : DFF_X1 port map( D => n2252, CK => CLK, Q => n9684
                           , QN => n14472);
   REGISTERS_reg_3_13_inst : DFF_X1 port map( D => n2251, CK => CLK, Q => n9683
                           , QN => n14471);
   REGISTERS_reg_3_12_inst : DFF_X1 port map( D => n2250, CK => CLK, Q => n9682
                           , QN => n14470);
   REGISTERS_reg_3_11_inst : DFF_X1 port map( D => n2249, CK => CLK, Q => n9681
                           , QN => n14469);
   REGISTERS_reg_3_10_inst : DFF_X1 port map( D => n2248, CK => CLK, Q => n9680
                           , QN => n14468);
   REGISTERS_reg_3_9_inst : DFF_X1 port map( D => n2247, CK => CLK, Q => n9679,
                           QN => n14467);
   REGISTERS_reg_3_8_inst : DFF_X1 port map( D => n2246, CK => CLK, Q => n9678,
                           QN => n14466);
   REGISTERS_reg_3_7_inst : DFF_X1 port map( D => n2245, CK => CLK, Q => n9677,
                           QN => n14465);
   REGISTERS_reg_3_6_inst : DFF_X1 port map( D => n2244, CK => CLK, Q => n9676,
                           QN => n14464);
   REGISTERS_reg_3_5_inst : DFF_X1 port map( D => n2243, CK => CLK, Q => n9675,
                           QN => n14463);
   REGISTERS_reg_3_4_inst : DFF_X1 port map( D => n2242, CK => CLK, Q => n9674,
                           QN => n14462);
   REGISTERS_reg_3_3_inst : DFF_X1 port map( D => n2241, CK => CLK, Q => n9673,
                           QN => n14461);
   REGISTERS_reg_3_2_inst : DFF_X1 port map( D => n2240, CK => CLK, Q => n9672,
                           QN => n14460);
   REGISTERS_reg_3_1_inst : DFF_X1 port map( D => n2239, CK => CLK, Q => n9671,
                           QN => n14459);
   REGISTERS_reg_3_0_inst : DFF_X1 port map( D => n2238, CK => CLK, Q => n9670,
                           QN => n14458);
   REGISTERS_reg_4_31_inst : DFF_X1 port map( D => n2237, CK => CLK, Q => 
                           n13323, QN => n14027);
   REGISTERS_reg_4_30_inst : DFF_X1 port map( D => n2236, CK => CLK, Q => 
                           n13322, QN => n14026);
   REGISTERS_reg_4_29_inst : DFF_X1 port map( D => n2235, CK => CLK, Q => 
                           n13321, QN => n14025);
   REGISTERS_reg_4_28_inst : DFF_X1 port map( D => n2234, CK => CLK, Q => 
                           n13320, QN => n14024);
   REGISTERS_reg_4_27_inst : DFF_X1 port map( D => n2233, CK => CLK, Q => 
                           n13319, QN => n14023);
   REGISTERS_reg_4_26_inst : DFF_X1 port map( D => n2232, CK => CLK, Q => 
                           n13318, QN => n14022);
   REGISTERS_reg_4_25_inst : DFF_X1 port map( D => n2231, CK => CLK, Q => 
                           n13317, QN => n14021);
   REGISTERS_reg_4_24_inst : DFF_X1 port map( D => n2230, CK => CLK, Q => 
                           n13316, QN => n14020);
   REGISTERS_reg_4_23_inst : DFF_X1 port map( D => n2229, CK => CLK, Q => 
                           n13419, QN => n14529);
   REGISTERS_reg_4_22_inst : DFF_X1 port map( D => n2228, CK => CLK, Q => 
                           n13418, QN => n14528);
   REGISTERS_reg_4_21_inst : DFF_X1 port map( D => n2227, CK => CLK, Q => 
                           n13417, QN => n14527);
   REGISTERS_reg_4_20_inst : DFF_X1 port map( D => n2226, CK => CLK, Q => 
                           n13416, QN => n14526);
   REGISTERS_reg_4_19_inst : DFF_X1 port map( D => n2225, CK => CLK, Q => 
                           n13415, QN => n14525);
   REGISTERS_reg_4_18_inst : DFF_X1 port map( D => n2224, CK => CLK, Q => 
                           n13414, QN => n14524);
   REGISTERS_reg_4_17_inst : DFF_X1 port map( D => n2223, CK => CLK, Q => 
                           n13413, QN => n14523);
   REGISTERS_reg_4_16_inst : DFF_X1 port map( D => n2222, CK => CLK, Q => 
                           n13412, QN => n14522);
   REGISTERS_reg_4_15_inst : DFF_X1 port map( D => n2221, CK => CLK, Q => 
                           n13411, QN => n14521);
   REGISTERS_reg_4_14_inst : DFF_X1 port map( D => n2220, CK => CLK, Q => 
                           n13410, QN => n14520);
   REGISTERS_reg_4_13_inst : DFF_X1 port map( D => n2219, CK => CLK, Q => 
                           n13409, QN => n14519);
   REGISTERS_reg_4_12_inst : DFF_X1 port map( D => n2218, CK => CLK, Q => 
                           n13408, QN => n14518);
   REGISTERS_reg_4_11_inst : DFF_X1 port map( D => n2217, CK => CLK, Q => 
                           n13407, QN => n14517);
   REGISTERS_reg_4_10_inst : DFF_X1 port map( D => n2216, CK => CLK, Q => 
                           n13406, QN => n14516);
   REGISTERS_reg_4_9_inst : DFF_X1 port map( D => n2215, CK => CLK, Q => n13405
                           , QN => n14515);
   REGISTERS_reg_4_8_inst : DFF_X1 port map( D => n2214, CK => CLK, Q => n13404
                           , QN => n14514);
   REGISTERS_reg_4_7_inst : DFF_X1 port map( D => n2213, CK => CLK, Q => n13403
                           , QN => n14513);
   REGISTERS_reg_4_6_inst : DFF_X1 port map( D => n2212, CK => CLK, Q => n13402
                           , QN => n14512);
   REGISTERS_reg_4_5_inst : DFF_X1 port map( D => n2211, CK => CLK, Q => n13401
                           , QN => n14511);
   REGISTERS_reg_4_4_inst : DFF_X1 port map( D => n2210, CK => CLK, Q => n13400
                           , QN => n14510);
   REGISTERS_reg_4_3_inst : DFF_X1 port map( D => n2209, CK => CLK, Q => n13399
                           , QN => n14509);
   REGISTERS_reg_4_2_inst : DFF_X1 port map( D => n2208, CK => CLK, Q => n13398
                           , QN => n14508);
   REGISTERS_reg_4_1_inst : DFF_X1 port map( D => n2207, CK => CLK, Q => n13397
                           , QN => n14507);
   REGISTERS_reg_4_0_inst : DFF_X1 port map( D => n2206, CK => CLK, Q => n13396
                           , QN => n14506);
   REGISTERS_reg_5_31_inst : DFF_X1 port map( D => n2205, CK => CLK, Q => 
                           n13315, QN => n13987);
   REGISTERS_reg_5_30_inst : DFF_X1 port map( D => n2204, CK => CLK, Q => 
                           n13314, QN => n13986);
   REGISTERS_reg_5_29_inst : DFF_X1 port map( D => n2203, CK => CLK, Q => 
                           n13313, QN => n13985);
   REGISTERS_reg_5_28_inst : DFF_X1 port map( D => n2202, CK => CLK, Q => 
                           n13312, QN => n13984);
   REGISTERS_reg_5_27_inst : DFF_X1 port map( D => n2201, CK => CLK, Q => 
                           n13311, QN => n13983);
   REGISTERS_reg_5_26_inst : DFF_X1 port map( D => n2200, CK => CLK, Q => 
                           n13310, QN => n13982);
   REGISTERS_reg_5_25_inst : DFF_X1 port map( D => n2199, CK => CLK, Q => 
                           n13309, QN => n13981);
   REGISTERS_reg_5_24_inst : DFF_X1 port map( D => n2198, CK => CLK, Q => 
                           n13308, QN => n13980);
   REGISTERS_reg_5_23_inst : DFF_X1 port map( D => n2197, CK => CLK, Q => 
                           n13395, QN => n14409);
   REGISTERS_reg_5_22_inst : DFF_X1 port map( D => n2196, CK => CLK, Q => 
                           n13394, QN => n14408);
   REGISTERS_reg_5_21_inst : DFF_X1 port map( D => n2195, CK => CLK, Q => 
                           n13393, QN => n14407);
   REGISTERS_reg_5_20_inst : DFF_X1 port map( D => n2194, CK => CLK, Q => 
                           n13392, QN => n14406);
   REGISTERS_reg_5_19_inst : DFF_X1 port map( D => n2193, CK => CLK, Q => 
                           n13391, QN => n14405);
   REGISTERS_reg_5_18_inst : DFF_X1 port map( D => n2192, CK => CLK, Q => 
                           n13390, QN => n14404);
   REGISTERS_reg_5_17_inst : DFF_X1 port map( D => n2191, CK => CLK, Q => 
                           n13389, QN => n14403);
   REGISTERS_reg_5_16_inst : DFF_X1 port map( D => n2190, CK => CLK, Q => 
                           n13388, QN => n14402);
   REGISTERS_reg_5_15_inst : DFF_X1 port map( D => n2189, CK => CLK, Q => 
                           n13387, QN => n14401);
   REGISTERS_reg_5_14_inst : DFF_X1 port map( D => n2188, CK => CLK, Q => 
                           n13386, QN => n14400);
   REGISTERS_reg_5_13_inst : DFF_X1 port map( D => n2187, CK => CLK, Q => 
                           n13385, QN => n14399);
   REGISTERS_reg_5_12_inst : DFF_X1 port map( D => n2186, CK => CLK, Q => 
                           n13384, QN => n14398);
   REGISTERS_reg_5_11_inst : DFF_X1 port map( D => n2185, CK => CLK, Q => 
                           n13383, QN => n14397);
   REGISTERS_reg_5_10_inst : DFF_X1 port map( D => n2184, CK => CLK, Q => 
                           n13382, QN => n14396);
   REGISTERS_reg_5_9_inst : DFF_X1 port map( D => n2183, CK => CLK, Q => n13381
                           , QN => n14395);
   REGISTERS_reg_5_8_inst : DFF_X1 port map( D => n2182, CK => CLK, Q => n13380
                           , QN => n14394);
   REGISTERS_reg_5_7_inst : DFF_X1 port map( D => n2181, CK => CLK, Q => n13379
                           , QN => n14393);
   REGISTERS_reg_5_6_inst : DFF_X1 port map( D => n2180, CK => CLK, Q => n13378
                           , QN => n14392);
   REGISTERS_reg_5_5_inst : DFF_X1 port map( D => n2179, CK => CLK, Q => n13377
                           , QN => n14391);
   REGISTERS_reg_5_4_inst : DFF_X1 port map( D => n2178, CK => CLK, Q => n13376
                           , QN => n14390);
   REGISTERS_reg_5_3_inst : DFF_X1 port map( D => n2177, CK => CLK, Q => n13375
                           , QN => n14389);
   REGISTERS_reg_5_2_inst : DFF_X1 port map( D => n2176, CK => CLK, Q => n13374
                           , QN => n14388);
   REGISTERS_reg_5_1_inst : DFF_X1 port map( D => n2175, CK => CLK, Q => n13373
                           , QN => n14387);
   REGISTERS_reg_5_0_inst : DFF_X1 port map( D => n2174, CK => CLK, Q => n13372
                           , QN => n14386);
   REGISTERS_reg_6_31_inst : DFF_X1 port map( D => n2173, CK => CLK, Q => 
                           n13307, QN => n14043);
   REGISTERS_reg_6_30_inst : DFF_X1 port map( D => n2172, CK => CLK, Q => 
                           n13306, QN => n14042);
   REGISTERS_reg_6_29_inst : DFF_X1 port map( D => n2171, CK => CLK, Q => 
                           n13305, QN => n14041);
   REGISTERS_reg_6_28_inst : DFF_X1 port map( D => n2170, CK => CLK, Q => 
                           n13304, QN => n14040);
   REGISTERS_reg_6_27_inst : DFF_X1 port map( D => n2169, CK => CLK, Q => 
                           n13303, QN => n14039);
   REGISTERS_reg_6_26_inst : DFF_X1 port map( D => n2168, CK => CLK, Q => 
                           n13302, QN => n14038);
   REGISTERS_reg_6_25_inst : DFF_X1 port map( D => n2167, CK => CLK, Q => 
                           n13301, QN => n14037);
   REGISTERS_reg_6_24_inst : DFF_X1 port map( D => n2166, CK => CLK, Q => 
                           n13300, QN => n14036);
   REGISTERS_reg_6_23_inst : DFF_X1 port map( D => n2165, CK => CLK, Q => 
                           n13371, QN => n14577);
   REGISTERS_reg_6_22_inst : DFF_X1 port map( D => n2164, CK => CLK, Q => 
                           n13370, QN => n14576);
   REGISTERS_reg_6_21_inst : DFF_X1 port map( D => n2163, CK => CLK, Q => 
                           n13369, QN => n14575);
   REGISTERS_reg_6_20_inst : DFF_X1 port map( D => n2162, CK => CLK, Q => 
                           n13368, QN => n14574);
   REGISTERS_reg_6_19_inst : DFF_X1 port map( D => n2161, CK => CLK, Q => 
                           n13367, QN => n14573);
   REGISTERS_reg_6_18_inst : DFF_X1 port map( D => n2160, CK => CLK, Q => 
                           n13366, QN => n14572);
   REGISTERS_reg_6_17_inst : DFF_X1 port map( D => n2159, CK => CLK, Q => 
                           n13365, QN => n14571);
   REGISTERS_reg_6_16_inst : DFF_X1 port map( D => n2158, CK => CLK, Q => 
                           n13364, QN => n14570);
   REGISTERS_reg_6_15_inst : DFF_X1 port map( D => n2157, CK => CLK, Q => 
                           n13363, QN => n14569);
   REGISTERS_reg_6_14_inst : DFF_X1 port map( D => n2156, CK => CLK, Q => 
                           n13362, QN => n14568);
   REGISTERS_reg_6_13_inst : DFF_X1 port map( D => n2155, CK => CLK, Q => 
                           n13361, QN => n14567);
   REGISTERS_reg_6_12_inst : DFF_X1 port map( D => n2154, CK => CLK, Q => 
                           n13360, QN => n14566);
   REGISTERS_reg_6_11_inst : DFF_X1 port map( D => n2153, CK => CLK, Q => 
                           n13359, QN => n14565);
   REGISTERS_reg_6_10_inst : DFF_X1 port map( D => n2152, CK => CLK, Q => 
                           n13358, QN => n14564);
   REGISTERS_reg_6_9_inst : DFF_X1 port map( D => n2151, CK => CLK, Q => n13357
                           , QN => n14563);
   REGISTERS_reg_6_8_inst : DFF_X1 port map( D => n2150, CK => CLK, Q => n13356
                           , QN => n14562);
   REGISTERS_reg_6_7_inst : DFF_X1 port map( D => n2149, CK => CLK, Q => n13355
                           , QN => n14561);
   REGISTERS_reg_6_6_inst : DFF_X1 port map( D => n2148, CK => CLK, Q => n13354
                           , QN => n14560);
   REGISTERS_reg_6_5_inst : DFF_X1 port map( D => n2147, CK => CLK, Q => n13353
                           , QN => n14559);
   REGISTERS_reg_6_4_inst : DFF_X1 port map( D => n2146, CK => CLK, Q => n13352
                           , QN => n14558);
   REGISTERS_reg_6_3_inst : DFF_X1 port map( D => n2145, CK => CLK, Q => n13351
                           , QN => n14557);
   REGISTERS_reg_6_2_inst : DFF_X1 port map( D => n2144, CK => CLK, Q => n13350
                           , QN => n14556);
   REGISTERS_reg_6_1_inst : DFF_X1 port map( D => n2143, CK => CLK, Q => n13349
                           , QN => n14555);
   REGISTERS_reg_6_0_inst : DFF_X1 port map( D => n2142, CK => CLK, Q => n13348
                           , QN => n14554);
   REGISTERS_reg_7_31_inst : DFF_X1 port map( D => n2141, CK => CLK, Q => n9895
                           , QN => n14003);
   REGISTERS_reg_7_30_inst : DFF_X1 port map( D => n2140, CK => CLK, Q => n9893
                           , QN => n14002);
   REGISTERS_reg_7_29_inst : DFF_X1 port map( D => n2139, CK => CLK, Q => n9955
                           , QN => n14001);
   REGISTERS_reg_7_28_inst : DFF_X1 port map( D => n2138, CK => CLK, Q => n9953
                           , QN => n14000);
   REGISTERS_reg_7_27_inst : DFF_X1 port map( D => n2137, CK => CLK, Q => n9951
                           , QN => n13999);
   REGISTERS_reg_7_26_inst : DFF_X1 port map( D => n2136, CK => CLK, Q => n9949
                           , QN => n13998);
   REGISTERS_reg_7_25_inst : DFF_X1 port map( D => n2135, CK => CLK, Q => n9947
                           , QN => n13997);
   REGISTERS_reg_7_24_inst : DFF_X1 port map( D => n2134, CK => CLK, Q => n9945
                           , QN => n13996);
   REGISTERS_reg_7_23_inst : DFF_X1 port map( D => n2133, CK => CLK, Q => n9943
                           , QN => n14457);
   REGISTERS_reg_7_22_inst : DFF_X1 port map( D => n2132, CK => CLK, Q => n9941
                           , QN => n14456);
   REGISTERS_reg_7_21_inst : DFF_X1 port map( D => n2131, CK => CLK, Q => n9939
                           , QN => n14455);
   REGISTERS_reg_7_20_inst : DFF_X1 port map( D => n2130, CK => CLK, Q => n9937
                           , QN => n14454);
   REGISTERS_reg_7_19_inst : DFF_X1 port map( D => n2129, CK => CLK, Q => n9935
                           , QN => n14453);
   REGISTERS_reg_7_18_inst : DFF_X1 port map( D => n2128, CK => CLK, Q => n9933
                           , QN => n14452);
   REGISTERS_reg_7_17_inst : DFF_X1 port map( D => n2127, CK => CLK, Q => n9931
                           , QN => n14451);
   REGISTERS_reg_7_16_inst : DFF_X1 port map( D => n2126, CK => CLK, Q => n9929
                           , QN => n14450);
   REGISTERS_reg_7_15_inst : DFF_X1 port map( D => n2125, CK => CLK, Q => n9927
                           , QN => n14449);
   REGISTERS_reg_7_14_inst : DFF_X1 port map( D => n2124, CK => CLK, Q => n9925
                           , QN => n14448);
   REGISTERS_reg_7_13_inst : DFF_X1 port map( D => n2123, CK => CLK, Q => n9923
                           , QN => n14447);
   REGISTERS_reg_7_12_inst : DFF_X1 port map( D => n2122, CK => CLK, Q => n9921
                           , QN => n14446);
   REGISTERS_reg_7_11_inst : DFF_X1 port map( D => n2121, CK => CLK, Q => n9919
                           , QN => n14445);
   REGISTERS_reg_7_10_inst : DFF_X1 port map( D => n2120, CK => CLK, Q => n9917
                           , QN => n14444);
   REGISTERS_reg_7_9_inst : DFF_X1 port map( D => n2119, CK => CLK, Q => n9915,
                           QN => n14443);
   REGISTERS_reg_7_8_inst : DFF_X1 port map( D => n2118, CK => CLK, Q => n9913,
                           QN => n14442);
   REGISTERS_reg_7_7_inst : DFF_X1 port map( D => n2117, CK => CLK, Q => n9911,
                           QN => n14441);
   REGISTERS_reg_7_6_inst : DFF_X1 port map( D => n2116, CK => CLK, Q => n9909,
                           QN => n14440);
   REGISTERS_reg_7_5_inst : DFF_X1 port map( D => n2115, CK => CLK, Q => n9907,
                           QN => n14439);
   REGISTERS_reg_7_4_inst : DFF_X1 port map( D => n2114, CK => CLK, Q => n9905,
                           QN => n14438);
   REGISTERS_reg_7_3_inst : DFF_X1 port map( D => n2113, CK => CLK, Q => n9903,
                           QN => n14437);
   REGISTERS_reg_7_2_inst : DFF_X1 port map( D => n2112, CK => CLK, Q => n9901,
                           QN => n14436);
   REGISTERS_reg_7_1_inst : DFF_X1 port map( D => n2111, CK => CLK, Q => n9899,
                           QN => n14435);
   REGISTERS_reg_7_0_inst : DFF_X1 port map( D => n2110, CK => CLK, Q => n9897,
                           QN => n14434);
   REGISTERS_reg_8_31_inst : DFF_X1 port map( D => n2109, CK => CLK, Q => 
                           n_1096, QN => n13759);
   REGISTERS_reg_8_30_inst : DFF_X1 port map( D => n2108, CK => CLK, Q => 
                           n_1097, QN => n13758);
   REGISTERS_reg_8_29_inst : DFF_X1 port map( D => n2107, CK => CLK, Q => 
                           n_1098, QN => n13757);
   REGISTERS_reg_8_28_inst : DFF_X1 port map( D => n2106, CK => CLK, Q => 
                           n_1099, QN => n13756);
   REGISTERS_reg_8_27_inst : DFF_X1 port map( D => n2105, CK => CLK, Q => 
                           n_1100, QN => n13755);
   REGISTERS_reg_8_26_inst : DFF_X1 port map( D => n2104, CK => CLK, Q => 
                           n_1101, QN => n13754);
   REGISTERS_reg_8_25_inst : DFF_X1 port map( D => n2103, CK => CLK, Q => 
                           n_1102, QN => n13753);
   REGISTERS_reg_8_24_inst : DFF_X1 port map( D => n2102, CK => CLK, Q => 
                           n_1103, QN => n13752);
   REGISTERS_reg_8_23_inst : DFF_X1 port map( D => n2101, CK => CLK, Q => 
                           n_1104, QN => n13779);
   REGISTERS_reg_8_22_inst : DFF_X1 port map( D => n2100, CK => CLK, Q => 
                           n_1105, QN => n13778);
   REGISTERS_reg_8_21_inst : DFF_X1 port map( D => n2099, CK => CLK, Q => 
                           n_1106, QN => n13777);
   REGISTERS_reg_8_20_inst : DFF_X1 port map( D => n2098, CK => CLK, Q => 
                           n_1107, QN => n13776);
   REGISTERS_reg_8_19_inst : DFF_X1 port map( D => n2097, CK => CLK, Q => 
                           n_1108, QN => n13775);
   REGISTERS_reg_8_18_inst : DFF_X1 port map( D => n2096, CK => CLK, Q => 
                           n_1109, QN => n13774);
   REGISTERS_reg_8_17_inst : DFF_X1 port map( D => n2095, CK => CLK, Q => 
                           n_1110, QN => n13773);
   REGISTERS_reg_8_16_inst : DFF_X1 port map( D => n2094, CK => CLK, Q => 
                           n_1111, QN => n13772);
   REGISTERS_reg_8_15_inst : DFF_X1 port map( D => n2093, CK => CLK, Q => 
                           n_1112, QN => n13771);
   REGISTERS_reg_8_14_inst : DFF_X1 port map( D => n2092, CK => CLK, Q => 
                           n_1113, QN => n13770);
   REGISTERS_reg_8_13_inst : DFF_X1 port map( D => n2091, CK => CLK, Q => 
                           n_1114, QN => n13769);
   REGISTERS_reg_8_12_inst : DFF_X1 port map( D => n2090, CK => CLK, Q => 
                           n_1115, QN => n13768);
   REGISTERS_reg_8_11_inst : DFF_X1 port map( D => n2089, CK => CLK, Q => 
                           n_1116, QN => n13843);
   REGISTERS_reg_8_10_inst : DFF_X1 port map( D => n2088, CK => CLK, Q => 
                           n_1117, QN => n13842);
   REGISTERS_reg_8_9_inst : DFF_X1 port map( D => n2087, CK => CLK, Q => n_1118
                           , QN => n13841);
   REGISTERS_reg_8_8_inst : DFF_X1 port map( D => n2086, CK => CLK, Q => n_1119
                           , QN => n13840);
   REGISTERS_reg_8_7_inst : DFF_X1 port map( D => n2085, CK => CLK, Q => n_1120
                           , QN => n13839);
   REGISTERS_reg_8_6_inst : DFF_X1 port map( D => n2084, CK => CLK, Q => n_1121
                           , QN => n13838);
   REGISTERS_reg_8_5_inst : DFF_X1 port map( D => n2083, CK => CLK, Q => n_1122
                           , QN => n13837);
   REGISTERS_reg_8_4_inst : DFF_X1 port map( D => n2082, CK => CLK, Q => n_1123
                           , QN => n13836);
   REGISTERS_reg_8_3_inst : DFF_X1 port map( D => n2081, CK => CLK, Q => n_1124
                           , QN => n13835);
   REGISTERS_reg_8_2_inst : DFF_X1 port map( D => n2080, CK => CLK, Q => n_1125
                           , QN => n13834);
   REGISTERS_reg_8_1_inst : DFF_X1 port map( D => n2079, CK => CLK, Q => n_1126
                           , QN => n13833);
   REGISTERS_reg_8_0_inst : DFF_X1 port map( D => n2078, CK => CLK, Q => n_1127
                           , QN => n13832);
   REGISTERS_reg_9_31_inst : DFF_X1 port map( D => n2077, CK => CLK, Q => 
                           n_1128, QN => n13863);
   REGISTERS_reg_9_30_inst : DFF_X1 port map( D => n2076, CK => CLK, Q => 
                           n_1129, QN => n13862);
   REGISTERS_reg_9_29_inst : DFF_X1 port map( D => n2075, CK => CLK, Q => 
                           n_1130, QN => n13861);
   REGISTERS_reg_9_28_inst : DFF_X1 port map( D => n2074, CK => CLK, Q => 
                           n_1131, QN => n13860);
   REGISTERS_reg_9_27_inst : DFF_X1 port map( D => n2073, CK => CLK, Q => 
                           n_1132, QN => n13859);
   REGISTERS_reg_9_26_inst : DFF_X1 port map( D => n2072, CK => CLK, Q => 
                           n_1133, QN => n13858);
   REGISTERS_reg_9_25_inst : DFF_X1 port map( D => n2071, CK => CLK, Q => 
                           n_1134, QN => n13857);
   REGISTERS_reg_9_24_inst : DFF_X1 port map( D => n2070, CK => CLK, Q => 
                           n_1135, QN => n13856);
   REGISTERS_reg_9_23_inst : DFF_X1 port map( D => n2069, CK => CLK, Q => 
                           n_1136, QN => n14117);
   REGISTERS_reg_9_22_inst : DFF_X1 port map( D => n2068, CK => CLK, Q => 
                           n_1137, QN => n14116);
   REGISTERS_reg_9_21_inst : DFF_X1 port map( D => n2067, CK => CLK, Q => 
                           n_1138, QN => n14115);
   REGISTERS_reg_9_20_inst : DFF_X1 port map( D => n2066, CK => CLK, Q => 
                           n_1139, QN => n14114);
   REGISTERS_reg_9_19_inst : DFF_X1 port map( D => n2065, CK => CLK, Q => 
                           n_1140, QN => n14113);
   REGISTERS_reg_9_18_inst : DFF_X1 port map( D => n2064, CK => CLK, Q => 
                           n_1141, QN => n14112);
   REGISTERS_reg_9_17_inst : DFF_X1 port map( D => n2063, CK => CLK, Q => 
                           n_1142, QN => n14111);
   REGISTERS_reg_9_16_inst : DFF_X1 port map( D => n2062, CK => CLK, Q => 
                           n_1143, QN => n14110);
   REGISTERS_reg_9_15_inst : DFF_X1 port map( D => n2061, CK => CLK, Q => 
                           n_1144, QN => n14109);
   REGISTERS_reg_9_14_inst : DFF_X1 port map( D => n2060, CK => CLK, Q => 
                           n_1145, QN => n14108);
   REGISTERS_reg_9_13_inst : DFF_X1 port map( D => n2059, CK => CLK, Q => 
                           n_1146, QN => n14107);
   REGISTERS_reg_9_12_inst : DFF_X1 port map( D => n2058, CK => CLK, Q => 
                           n_1147, QN => n14106);
   REGISTERS_reg_9_11_inst : DFF_X1 port map( D => n2057, CK => CLK, Q => 
                           n_1148, QN => n14105);
   REGISTERS_reg_9_10_inst : DFF_X1 port map( D => n2056, CK => CLK, Q => 
                           n_1149, QN => n14104);
   REGISTERS_reg_9_9_inst : DFF_X1 port map( D => n2055, CK => CLK, Q => n_1150
                           , QN => n14103);
   REGISTERS_reg_9_8_inst : DFF_X1 port map( D => n2054, CK => CLK, Q => n_1151
                           , QN => n14102);
   REGISTERS_reg_9_7_inst : DFF_X1 port map( D => n2053, CK => CLK, Q => n_1152
                           , QN => n14101);
   REGISTERS_reg_9_6_inst : DFF_X1 port map( D => n2052, CK => CLK, Q => n_1153
                           , QN => n14100);
   REGISTERS_reg_9_5_inst : DFF_X1 port map( D => n2051, CK => CLK, Q => n_1154
                           , QN => n14099);
   REGISTERS_reg_9_4_inst : DFF_X1 port map( D => n2050, CK => CLK, Q => n_1155
                           , QN => n14098);
   REGISTERS_reg_9_3_inst : DFF_X1 port map( D => n2049, CK => CLK, Q => n_1156
                           , QN => n14097);
   REGISTERS_reg_9_2_inst : DFF_X1 port map( D => n2048, CK => CLK, Q => n_1157
                           , QN => n14096);
   REGISTERS_reg_9_1_inst : DFF_X1 port map( D => n2047, CK => CLK, Q => n_1158
                           , QN => n14095);
   REGISTERS_reg_9_0_inst : DFF_X1 port map( D => n2046, CK => CLK, Q => n_1159
                           , QN => n14094);
   REGISTERS_reg_10_31_inst : DFF_X1 port map( D => n2045, CK => CLK, Q => 
                           n_1160, QN => n13659);
   REGISTERS_reg_10_30_inst : DFF_X1 port map( D => n2044, CK => CLK, Q => 
                           n_1161, QN => n13658);
   REGISTERS_reg_10_29_inst : DFF_X1 port map( D => n2043, CK => CLK, Q => 
                           n_1162, QN => n13657);
   REGISTERS_reg_10_28_inst : DFF_X1 port map( D => n2042, CK => CLK, Q => 
                           n_1163, QN => n13656);
   REGISTERS_reg_10_27_inst : DFF_X1 port map( D => n2041, CK => CLK, Q => 
                           n_1164, QN => n13655);
   REGISTERS_reg_10_26_inst : DFF_X1 port map( D => n2040, CK => CLK, Q => 
                           n_1165, QN => n13654);
   REGISTERS_reg_10_25_inst : DFF_X1 port map( D => n2039, CK => CLK, Q => 
                           n_1166, QN => n13653);
   REGISTERS_reg_10_24_inst : DFF_X1 port map( D => n2038, CK => CLK, Q => 
                           n_1167, QN => n13652);
   REGISTERS_reg_10_23_inst : DFF_X1 port map( D => n2037, CK => CLK, Q => 
                           n_1168, QN => n13683);
   REGISTERS_reg_10_22_inst : DFF_X1 port map( D => n2036, CK => CLK, Q => 
                           n_1169, QN => n13682);
   REGISTERS_reg_10_21_inst : DFF_X1 port map( D => n2035, CK => CLK, Q => 
                           n_1170, QN => n13681);
   REGISTERS_reg_10_20_inst : DFF_X1 port map( D => n2034, CK => CLK, Q => 
                           n_1171, QN => n13680);
   REGISTERS_reg_10_19_inst : DFF_X1 port map( D => n2033, CK => CLK, Q => 
                           n_1172, QN => n13679);
   REGISTERS_reg_10_18_inst : DFF_X1 port map( D => n2032, CK => CLK, Q => 
                           n_1173, QN => n13678);
   REGISTERS_reg_10_17_inst : DFF_X1 port map( D => n2031, CK => CLK, Q => 
                           n_1174, QN => n13677);
   REGISTERS_reg_10_16_inst : DFF_X1 port map( D => n2030, CK => CLK, Q => 
                           n_1175, QN => n13676);
   REGISTERS_reg_10_15_inst : DFF_X1 port map( D => n2029, CK => CLK, Q => 
                           n_1176, QN => n13675);
   REGISTERS_reg_10_14_inst : DFF_X1 port map( D => n2028, CK => CLK, Q => 
                           n_1177, QN => n13674);
   REGISTERS_reg_10_13_inst : DFF_X1 port map( D => n2027, CK => CLK, Q => 
                           n_1178, QN => n13673);
   REGISTERS_reg_10_12_inst : DFF_X1 port map( D => n2026, CK => CLK, Q => 
                           n_1179, QN => n13672);
   REGISTERS_reg_10_11_inst : DFF_X1 port map( D => n2025, CK => CLK, Q => 
                           n_1180, QN => n13751);
   REGISTERS_reg_10_10_inst : DFF_X1 port map( D => n2024, CK => CLK, Q => 
                           n_1181, QN => n13750);
   REGISTERS_reg_10_9_inst : DFF_X1 port map( D => n2023, CK => CLK, Q => 
                           n_1182, QN => n13749);
   REGISTERS_reg_10_8_inst : DFF_X1 port map( D => n2022, CK => CLK, Q => 
                           n_1183, QN => n13748);
   REGISTERS_reg_10_7_inst : DFF_X1 port map( D => n2021, CK => CLK, Q => 
                           n_1184, QN => n13747);
   REGISTERS_reg_10_6_inst : DFF_X1 port map( D => n2020, CK => CLK, Q => 
                           n_1185, QN => n13746);
   REGISTERS_reg_10_5_inst : DFF_X1 port map( D => n2019, CK => CLK, Q => 
                           n_1186, QN => n13745);
   REGISTERS_reg_10_4_inst : DFF_X1 port map( D => n2018, CK => CLK, Q => 
                           n_1187, QN => n13744);
   REGISTERS_reg_10_3_inst : DFF_X1 port map( D => n2017, CK => CLK, Q => 
                           n_1188, QN => n13743);
   REGISTERS_reg_10_2_inst : DFF_X1 port map( D => n2016, CK => CLK, Q => 
                           n_1189, QN => n13742);
   REGISTERS_reg_10_1_inst : DFF_X1 port map( D => n2015, CK => CLK, Q => 
                           n_1190, QN => n13741);
   REGISTERS_reg_10_0_inst : DFF_X1 port map( D => n2014, CK => CLK, Q => 
                           n_1191, QN => n13740);
   REGISTERS_reg_11_31_inst : DFF_X1 port map( D => n2013, CK => CLK, Q => 
                           n14320, QN => n8988);
   REGISTERS_reg_11_30_inst : DFF_X1 port map( D => n2012, CK => CLK, Q => 
                           n14318, QN => n8989);
   REGISTERS_reg_11_29_inst : DFF_X1 port map( D => n2011, CK => CLK, Q => 
                           n14316, QN => n8990);
   REGISTERS_reg_11_28_inst : DFF_X1 port map( D => n2010, CK => CLK, Q => 
                           n14314, QN => n8991);
   REGISTERS_reg_11_27_inst : DFF_X1 port map( D => n2009, CK => CLK, Q => 
                           n14312, QN => n8992);
   REGISTERS_reg_11_26_inst : DFF_X1 port map( D => n2008, CK => CLK, Q => 
                           n14310, QN => n8993);
   REGISTERS_reg_11_25_inst : DFF_X1 port map( D => n2007, CK => CLK, Q => 
                           n14308, QN => n8994);
   REGISTERS_reg_11_24_inst : DFF_X1 port map( D => n2006, CK => CLK, Q => 
                           n14306, QN => n8995);
   REGISTERS_reg_11_23_inst : DFF_X1 port map( D => n2005, CK => CLK, Q => 
                           n14304, QN => n8996);
   REGISTERS_reg_11_22_inst : DFF_X1 port map( D => n2004, CK => CLK, Q => 
                           n14302, QN => n8997);
   REGISTERS_reg_11_21_inst : DFF_X1 port map( D => n2003, CK => CLK, Q => 
                           n14300, QN => n8998);
   REGISTERS_reg_11_20_inst : DFF_X1 port map( D => n2002, CK => CLK, Q => 
                           n14298, QN => n8999);
   REGISTERS_reg_11_19_inst : DFF_X1 port map( D => n2001, CK => CLK, Q => 
                           n14296, QN => n9000);
   REGISTERS_reg_11_18_inst : DFF_X1 port map( D => n2000, CK => CLK, Q => 
                           n14294, QN => n9001);
   REGISTERS_reg_11_17_inst : DFF_X1 port map( D => n1999, CK => CLK, Q => 
                           n14292, QN => n9002);
   REGISTERS_reg_11_16_inst : DFF_X1 port map( D => n1998, CK => CLK, Q => 
                           n14290, QN => n9003);
   REGISTERS_reg_11_15_inst : DFF_X1 port map( D => n1997, CK => CLK, Q => 
                           n14288, QN => n9004);
   REGISTERS_reg_11_14_inst : DFF_X1 port map( D => n1996, CK => CLK, Q => 
                           n14286, QN => n9005);
   REGISTERS_reg_11_13_inst : DFF_X1 port map( D => n1995, CK => CLK, Q => 
                           n14284, QN => n9006);
   REGISTERS_reg_11_12_inst : DFF_X1 port map( D => n1994, CK => CLK, Q => 
                           n14282, QN => n9007);
   REGISTERS_reg_11_11_inst : DFF_X1 port map( D => n1993, CK => CLK, Q => 
                           n14280, QN => n9008);
   REGISTERS_reg_11_10_inst : DFF_X1 port map( D => n1992, CK => CLK, Q => 
                           n14278, QN => n9009);
   REGISTERS_reg_11_9_inst : DFF_X1 port map( D => n1991, CK => CLK, Q => 
                           n14276, QN => n9010);
   REGISTERS_reg_11_8_inst : DFF_X1 port map( D => n1990, CK => CLK, Q => 
                           n14274, QN => n9011);
   REGISTERS_reg_11_7_inst : DFF_X1 port map( D => n1989, CK => CLK, Q => 
                           n14272, QN => n9012);
   REGISTERS_reg_11_6_inst : DFF_X1 port map( D => n1988, CK => CLK, Q => 
                           n14270, QN => n9013);
   REGISTERS_reg_11_5_inst : DFF_X1 port map( D => n1987, CK => CLK, Q => 
                           n14268, QN => n9014);
   REGISTERS_reg_11_4_inst : DFF_X1 port map( D => n1986, CK => CLK, Q => 
                           n14266, QN => n9015);
   REGISTERS_reg_11_3_inst : DFF_X1 port map( D => n1985, CK => CLK, Q => 
                           n14264, QN => n9016);
   REGISTERS_reg_11_2_inst : DFF_X1 port map( D => n1984, CK => CLK, Q => 
                           n14262, QN => n9017);
   REGISTERS_reg_11_1_inst : DFF_X1 port map( D => n1983, CK => CLK, Q => 
                           n14260, QN => n9018);
   REGISTERS_reg_11_0_inst : DFF_X1 port map( D => n1982, CK => CLK, Q => 
                           n14258, QN => n9019);
   REGISTERS_reg_12_31_inst : DFF_X1 port map( D => n1981, CK => CLK, Q => 
                           n13275, QN => n14019);
   REGISTERS_reg_12_30_inst : DFF_X1 port map( D => n1980, CK => CLK, Q => 
                           n13274, QN => n14018);
   REGISTERS_reg_12_29_inst : DFF_X1 port map( D => n1979, CK => CLK, Q => 
                           n13273, QN => n14017);
   REGISTERS_reg_12_28_inst : DFF_X1 port map( D => n1978, CK => CLK, Q => 
                           n13272, QN => n14016);
   REGISTERS_reg_12_27_inst : DFF_X1 port map( D => n1977, CK => CLK, Q => 
                           n13271, QN => n14015);
   REGISTERS_reg_12_26_inst : DFF_X1 port map( D => n1976, CK => CLK, Q => 
                           n13270, QN => n14014);
   REGISTERS_reg_12_25_inst : DFF_X1 port map( D => n1975, CK => CLK, Q => 
                           n13269, QN => n14013);
   REGISTERS_reg_12_24_inst : DFF_X1 port map( D => n1974, CK => CLK, Q => 
                           n13268, QN => n14012);
   REGISTERS_reg_12_23_inst : DFF_X1 port map( D => n1973, CK => CLK, Q => 
                           n13563, QN => n14505);
   REGISTERS_reg_12_22_inst : DFF_X1 port map( D => n1972, CK => CLK, Q => 
                           n13562, QN => n14504);
   REGISTERS_reg_12_21_inst : DFF_X1 port map( D => n1971, CK => CLK, Q => 
                           n13561, QN => n14503);
   REGISTERS_reg_12_20_inst : DFF_X1 port map( D => n1970, CK => CLK, Q => 
                           n13560, QN => n14502);
   REGISTERS_reg_12_19_inst : DFF_X1 port map( D => n1969, CK => CLK, Q => 
                           n13559, QN => n14501);
   REGISTERS_reg_12_18_inst : DFF_X1 port map( D => n1968, CK => CLK, Q => 
                           n13558, QN => n14500);
   REGISTERS_reg_12_17_inst : DFF_X1 port map( D => n1967, CK => CLK, Q => 
                           n13557, QN => n14499);
   REGISTERS_reg_12_16_inst : DFF_X1 port map( D => n1966, CK => CLK, Q => 
                           n13556, QN => n14498);
   REGISTERS_reg_12_15_inst : DFF_X1 port map( D => n1965, CK => CLK, Q => 
                           n13555, QN => n14497);
   REGISTERS_reg_12_14_inst : DFF_X1 port map( D => n1964, CK => CLK, Q => 
                           n13554, QN => n14496);
   REGISTERS_reg_12_13_inst : DFF_X1 port map( D => n1963, CK => CLK, Q => 
                           n13553, QN => n14495);
   REGISTERS_reg_12_12_inst : DFF_X1 port map( D => n1962, CK => CLK, Q => 
                           n13552, QN => n14494);
   REGISTERS_reg_12_11_inst : DFF_X1 port map( D => n1961, CK => CLK, Q => 
                           n13551, QN => n14493);
   REGISTERS_reg_12_10_inst : DFF_X1 port map( D => n1960, CK => CLK, Q => 
                           n13550, QN => n14492);
   REGISTERS_reg_12_9_inst : DFF_X1 port map( D => n1959, CK => CLK, Q => 
                           n13549, QN => n14491);
   REGISTERS_reg_12_8_inst : DFF_X1 port map( D => n1958, CK => CLK, Q => 
                           n13548, QN => n14490);
   REGISTERS_reg_12_7_inst : DFF_X1 port map( D => n1957, CK => CLK, Q => 
                           n13547, QN => n14489);
   REGISTERS_reg_12_6_inst : DFF_X1 port map( D => n1956, CK => CLK, Q => 
                           n13546, QN => n14488);
   REGISTERS_reg_12_5_inst : DFF_X1 port map( D => n1955, CK => CLK, Q => 
                           n13545, QN => n14487);
   REGISTERS_reg_12_4_inst : DFF_X1 port map( D => n1954, CK => CLK, Q => 
                           n13544, QN => n14486);
   REGISTERS_reg_12_3_inst : DFF_X1 port map( D => n1953, CK => CLK, Q => 
                           n13543, QN => n14485);
   REGISTERS_reg_12_2_inst : DFF_X1 port map( D => n1952, CK => CLK, Q => 
                           n13542, QN => n14484);
   REGISTERS_reg_12_1_inst : DFF_X1 port map( D => n1951, CK => CLK, Q => 
                           n13541, QN => n14483);
   REGISTERS_reg_12_0_inst : DFF_X1 port map( D => n1950, CK => CLK, Q => 
                           n13540, QN => n14482);
   REGISTERS_reg_13_31_inst : DFF_X1 port map( D => n1949, CK => CLK, Q => 
                           n13267, QN => n13995);
   REGISTERS_reg_13_30_inst : DFF_X1 port map( D => n1948, CK => CLK, Q => 
                           n13266, QN => n13994);
   REGISTERS_reg_13_29_inst : DFF_X1 port map( D => n1947, CK => CLK, Q => 
                           n13265, QN => n13993);
   REGISTERS_reg_13_28_inst : DFF_X1 port map( D => n1946, CK => CLK, Q => 
                           n13264, QN => n13992);
   REGISTERS_reg_13_27_inst : DFF_X1 port map( D => n1945, CK => CLK, Q => 
                           n13263, QN => n13991);
   REGISTERS_reg_13_26_inst : DFF_X1 port map( D => n1944, CK => CLK, Q => 
                           n13262, QN => n13990);
   REGISTERS_reg_13_25_inst : DFF_X1 port map( D => n1943, CK => CLK, Q => 
                           n13261, QN => n13989);
   REGISTERS_reg_13_24_inst : DFF_X1 port map( D => n1942, CK => CLK, Q => 
                           n13260, QN => n13988);
   REGISTERS_reg_13_23_inst : DFF_X1 port map( D => n1941, CK => CLK, Q => 
                           n13539, QN => n14433);
   REGISTERS_reg_13_22_inst : DFF_X1 port map( D => n1940, CK => CLK, Q => 
                           n13538, QN => n14432);
   REGISTERS_reg_13_21_inst : DFF_X1 port map( D => n1939, CK => CLK, Q => 
                           n13537, QN => n14431);
   REGISTERS_reg_13_20_inst : DFF_X1 port map( D => n1938, CK => CLK, Q => 
                           n13536, QN => n14430);
   REGISTERS_reg_13_19_inst : DFF_X1 port map( D => n1937, CK => CLK, Q => 
                           n13535, QN => n14429);
   REGISTERS_reg_13_18_inst : DFF_X1 port map( D => n1936, CK => CLK, Q => 
                           n13534, QN => n14428);
   REGISTERS_reg_13_17_inst : DFF_X1 port map( D => n1935, CK => CLK, Q => 
                           n13533, QN => n14427);
   REGISTERS_reg_13_16_inst : DFF_X1 port map( D => n1934, CK => CLK, Q => 
                           n13532, QN => n14426);
   REGISTERS_reg_13_15_inst : DFF_X1 port map( D => n1933, CK => CLK, Q => 
                           n13531, QN => n14425);
   REGISTERS_reg_13_14_inst : DFF_X1 port map( D => n1932, CK => CLK, Q => 
                           n13530, QN => n14424);
   REGISTERS_reg_13_13_inst : DFF_X1 port map( D => n1931, CK => CLK, Q => 
                           n13529, QN => n14423);
   REGISTERS_reg_13_12_inst : DFF_X1 port map( D => n1930, CK => CLK, Q => 
                           n13528, QN => n14422);
   REGISTERS_reg_13_11_inst : DFF_X1 port map( D => n1929, CK => CLK, Q => 
                           n13527, QN => n14421);
   REGISTERS_reg_13_10_inst : DFF_X1 port map( D => n1928, CK => CLK, Q => 
                           n13526, QN => n14420);
   REGISTERS_reg_13_9_inst : DFF_X1 port map( D => n1927, CK => CLK, Q => 
                           n13525, QN => n14419);
   REGISTERS_reg_13_8_inst : DFF_X1 port map( D => n1926, CK => CLK, Q => 
                           n13524, QN => n14418);
   REGISTERS_reg_13_7_inst : DFF_X1 port map( D => n1925, CK => CLK, Q => 
                           n13523, QN => n14417);
   REGISTERS_reg_13_6_inst : DFF_X1 port map( D => n1924, CK => CLK, Q => 
                           n13522, QN => n14416);
   REGISTERS_reg_13_5_inst : DFF_X1 port map( D => n1923, CK => CLK, Q => 
                           n13521, QN => n14415);
   REGISTERS_reg_13_4_inst : DFF_X1 port map( D => n1922, CK => CLK, Q => 
                           n13520, QN => n14414);
   REGISTERS_reg_13_3_inst : DFF_X1 port map( D => n1921, CK => CLK, Q => 
                           n13519, QN => n14413);
   REGISTERS_reg_13_2_inst : DFF_X1 port map( D => n1920, CK => CLK, Q => 
                           n13518, QN => n14412);
   REGISTERS_reg_13_1_inst : DFF_X1 port map( D => n1919, CK => CLK, Q => 
                           n13517, QN => n14411);
   REGISTERS_reg_13_0_inst : DFF_X1 port map( D => n1918, CK => CLK, Q => 
                           n13516, QN => n14410);
   REGISTERS_reg_14_31_inst : DFF_X1 port map( D => n1917, CK => CLK, Q => 
                           n13259, QN => n14035);
   REGISTERS_reg_14_30_inst : DFF_X1 port map( D => n1916, CK => CLK, Q => 
                           n13258, QN => n14034);
   REGISTERS_reg_14_29_inst : DFF_X1 port map( D => n1915, CK => CLK, Q => 
                           n13257, QN => n14033);
   REGISTERS_reg_14_28_inst : DFF_X1 port map( D => n1914, CK => CLK, Q => 
                           n13256, QN => n14032);
   REGISTERS_reg_14_27_inst : DFF_X1 port map( D => n1913, CK => CLK, Q => 
                           n13255, QN => n14031);
   REGISTERS_reg_14_26_inst : DFF_X1 port map( D => n1912, CK => CLK, Q => 
                           n13254, QN => n14030);
   REGISTERS_reg_14_25_inst : DFF_X1 port map( D => n1911, CK => CLK, Q => 
                           n13253, QN => n14029);
   REGISTERS_reg_14_24_inst : DFF_X1 port map( D => n1910, CK => CLK, Q => 
                           n13252, QN => n14028);
   REGISTERS_reg_14_23_inst : DFF_X1 port map( D => n1909, CK => CLK, Q => 
                           n13515, QN => n14553);
   REGISTERS_reg_14_22_inst : DFF_X1 port map( D => n1908, CK => CLK, Q => 
                           n13514, QN => n14552);
   REGISTERS_reg_14_21_inst : DFF_X1 port map( D => n1907, CK => CLK, Q => 
                           n13513, QN => n14551);
   REGISTERS_reg_14_20_inst : DFF_X1 port map( D => n1906, CK => CLK, Q => 
                           n13512, QN => n14550);
   REGISTERS_reg_14_19_inst : DFF_X1 port map( D => n1905, CK => CLK, Q => 
                           n13511, QN => n14549);
   REGISTERS_reg_14_18_inst : DFF_X1 port map( D => n1904, CK => CLK, Q => 
                           n13510, QN => n14548);
   REGISTERS_reg_14_17_inst : DFF_X1 port map( D => n1903, CK => CLK, Q => 
                           n13509, QN => n14547);
   REGISTERS_reg_14_16_inst : DFF_X1 port map( D => n1902, CK => CLK, Q => 
                           n13508, QN => n14546);
   REGISTERS_reg_14_15_inst : DFF_X1 port map( D => n1901, CK => CLK, Q => 
                           n13507, QN => n14545);
   REGISTERS_reg_14_14_inst : DFF_X1 port map( D => n1900, CK => CLK, Q => 
                           n13506, QN => n14544);
   REGISTERS_reg_14_13_inst : DFF_X1 port map( D => n1899, CK => CLK, Q => 
                           n13505, QN => n14543);
   REGISTERS_reg_14_12_inst : DFF_X1 port map( D => n1898, CK => CLK, Q => 
                           n13504, QN => n14542);
   REGISTERS_reg_14_11_inst : DFF_X1 port map( D => n1897, CK => CLK, Q => 
                           n13503, QN => n14541);
   REGISTERS_reg_14_10_inst : DFF_X1 port map( D => n1896, CK => CLK, Q => 
                           n13502, QN => n14540);
   REGISTERS_reg_14_9_inst : DFF_X1 port map( D => n1895, CK => CLK, Q => 
                           n13501, QN => n14539);
   REGISTERS_reg_14_8_inst : DFF_X1 port map( D => n1894, CK => CLK, Q => 
                           n13500, QN => n14538);
   REGISTERS_reg_14_7_inst : DFF_X1 port map( D => n1893, CK => CLK, Q => 
                           n13499, QN => n14537);
   REGISTERS_reg_14_6_inst : DFF_X1 port map( D => n1892, CK => CLK, Q => 
                           n13498, QN => n14536);
   REGISTERS_reg_14_5_inst : DFF_X1 port map( D => n1891, CK => CLK, Q => 
                           n13497, QN => n14535);
   REGISTERS_reg_14_4_inst : DFF_X1 port map( D => n1890, CK => CLK, Q => 
                           n13496, QN => n14534);
   REGISTERS_reg_14_3_inst : DFF_X1 port map( D => n1889, CK => CLK, Q => 
                           n13495, QN => n14533);
   REGISTERS_reg_14_2_inst : DFF_X1 port map( D => n1888, CK => CLK, Q => 
                           n13494, QN => n14532);
   REGISTERS_reg_14_1_inst : DFF_X1 port map( D => n1887, CK => CLK, Q => 
                           n13493, QN => n14531);
   REGISTERS_reg_14_0_inst : DFF_X1 port map( D => n1886, CK => CLK, Q => 
                           n13492, QN => n14530);
   REGISTERS_reg_15_31_inst : DFF_X1 port map( D => n1885, CK => CLK, Q => 
                           n14321, QN => n9116);
   REGISTERS_reg_15_30_inst : DFF_X1 port map( D => n1884, CK => CLK, Q => 
                           n14319, QN => n9117);
   REGISTERS_reg_15_29_inst : DFF_X1 port map( D => n1883, CK => CLK, Q => 
                           n14317, QN => n9118);
   REGISTERS_reg_15_28_inst : DFF_X1 port map( D => n1882, CK => CLK, Q => 
                           n14315, QN => n9119);
   REGISTERS_reg_15_27_inst : DFF_X1 port map( D => n1881, CK => CLK, Q => 
                           n14313, QN => n9120);
   REGISTERS_reg_15_26_inst : DFF_X1 port map( D => n1880, CK => CLK, Q => 
                           n14311, QN => n9121);
   REGISTERS_reg_15_25_inst : DFF_X1 port map( D => n1879, CK => CLK, Q => 
                           n14309, QN => n9122);
   REGISTERS_reg_15_24_inst : DFF_X1 port map( D => n1878, CK => CLK, Q => 
                           n14307, QN => n9123);
   REGISTERS_reg_15_23_inst : DFF_X1 port map( D => n1877, CK => CLK, Q => 
                           n14305, QN => n9124);
   REGISTERS_reg_15_22_inst : DFF_X1 port map( D => n1876, CK => CLK, Q => 
                           n14303, QN => n9125);
   REGISTERS_reg_15_21_inst : DFF_X1 port map( D => n1875, CK => CLK, Q => 
                           n14301, QN => n9126);
   REGISTERS_reg_15_20_inst : DFF_X1 port map( D => n1874, CK => CLK, Q => 
                           n14299, QN => n9127);
   REGISTERS_reg_15_19_inst : DFF_X1 port map( D => n1873, CK => CLK, Q => 
                           n14297, QN => n9128);
   REGISTERS_reg_15_18_inst : DFF_X1 port map( D => n1872, CK => CLK, Q => 
                           n14295, QN => n9129);
   REGISTERS_reg_15_17_inst : DFF_X1 port map( D => n1871, CK => CLK, Q => 
                           n14293, QN => n9130);
   REGISTERS_reg_15_16_inst : DFF_X1 port map( D => n1870, CK => CLK, Q => 
                           n14291, QN => n9131);
   REGISTERS_reg_15_15_inst : DFF_X1 port map( D => n1869, CK => CLK, Q => 
                           n14289, QN => n9132);
   REGISTERS_reg_15_14_inst : DFF_X1 port map( D => n1868, CK => CLK, Q => 
                           n14287, QN => n9133);
   REGISTERS_reg_15_13_inst : DFF_X1 port map( D => n1867, CK => CLK, Q => 
                           n14285, QN => n9134);
   REGISTERS_reg_15_12_inst : DFF_X1 port map( D => n1866, CK => CLK, Q => 
                           n14283, QN => n9135);
   REGISTERS_reg_15_11_inst : DFF_X1 port map( D => n1865, CK => CLK, Q => 
                           n14281, QN => n9136);
   REGISTERS_reg_15_10_inst : DFF_X1 port map( D => n1864, CK => CLK, Q => 
                           n14279, QN => n9137);
   REGISTERS_reg_15_9_inst : DFF_X1 port map( D => n1863, CK => CLK, Q => 
                           n14277, QN => n9138);
   REGISTERS_reg_15_8_inst : DFF_X1 port map( D => n1862, CK => CLK, Q => 
                           n14275, QN => n9139);
   REGISTERS_reg_15_7_inst : DFF_X1 port map( D => n1861, CK => CLK, Q => 
                           n14273, QN => n9140);
   REGISTERS_reg_15_6_inst : DFF_X1 port map( D => n1860, CK => CLK, Q => 
                           n14271, QN => n9141);
   REGISTERS_reg_15_5_inst : DFF_X1 port map( D => n1859, CK => CLK, Q => 
                           n14269, QN => n9142);
   REGISTERS_reg_15_4_inst : DFF_X1 port map( D => n1858, CK => CLK, Q => 
                           n14267, QN => n9143);
   REGISTERS_reg_15_3_inst : DFF_X1 port map( D => n1857, CK => CLK, Q => 
                           n14265, QN => n9144);
   REGISTERS_reg_15_2_inst : DFF_X1 port map( D => n1856, CK => CLK, Q => 
                           n14263, QN => n9145);
   REGISTERS_reg_15_1_inst : DFF_X1 port map( D => n1855, CK => CLK, Q => 
                           n14261, QN => n9146);
   REGISTERS_reg_15_0_inst : DFF_X1 port map( D => n1854, CK => CLK, Q => 
                           n14259, QN => n9147);
   REGISTERS_reg_16_31_inst : DFF_X1 port map( D => n1853, CK => CLK, Q => 
                           n_1192, QN => n13879);
   REGISTERS_reg_16_30_inst : DFF_X1 port map( D => n1852, CK => CLK, Q => 
                           n_1193, QN => n13878);
   REGISTERS_reg_16_29_inst : DFF_X1 port map( D => n1851, CK => CLK, Q => 
                           n_1194, QN => n13877);
   REGISTERS_reg_16_28_inst : DFF_X1 port map( D => n1850, CK => CLK, Q => 
                           n_1195, QN => n13876);
   REGISTERS_reg_16_27_inst : DFF_X1 port map( D => n1849, CK => CLK, Q => 
                           n_1196, QN => n13875);
   REGISTERS_reg_16_26_inst : DFF_X1 port map( D => n1848, CK => CLK, Q => 
                           n_1197, QN => n13874);
   REGISTERS_reg_16_25_inst : DFF_X1 port map( D => n1847, CK => CLK, Q => 
                           n_1198, QN => n13873);
   REGISTERS_reg_16_24_inst : DFF_X1 port map( D => n1846, CK => CLK, Q => 
                           n_1199, QN => n13872);
   REGISTERS_reg_16_23_inst : DFF_X1 port map( D => n1845, CK => CLK, Q => 
                           n_1200, QN => n14165);
   REGISTERS_reg_16_22_inst : DFF_X1 port map( D => n1844, CK => CLK, Q => 
                           n_1201, QN => n14164);
   REGISTERS_reg_16_21_inst : DFF_X1 port map( D => n1843, CK => CLK, Q => 
                           n_1202, QN => n14163);
   REGISTERS_reg_16_20_inst : DFF_X1 port map( D => n1842, CK => CLK, Q => 
                           n_1203, QN => n14162);
   REGISTERS_reg_16_19_inst : DFF_X1 port map( D => n1841, CK => CLK, Q => 
                           n_1204, QN => n14161);
   REGISTERS_reg_16_18_inst : DFF_X1 port map( D => n1840, CK => CLK, Q => 
                           n_1205, QN => n14160);
   REGISTERS_reg_16_17_inst : DFF_X1 port map( D => n1839, CK => CLK, Q => 
                           n_1206, QN => n14159);
   REGISTERS_reg_16_16_inst : DFF_X1 port map( D => n1838, CK => CLK, Q => 
                           n_1207, QN => n14158);
   REGISTERS_reg_16_15_inst : DFF_X1 port map( D => n1837, CK => CLK, Q => 
                           n_1208, QN => n14157);
   REGISTERS_reg_16_14_inst : DFF_X1 port map( D => n1836, CK => CLK, Q => 
                           n_1209, QN => n14156);
   REGISTERS_reg_16_13_inst : DFF_X1 port map( D => n1835, CK => CLK, Q => 
                           n_1210, QN => n14155);
   REGISTERS_reg_16_12_inst : DFF_X1 port map( D => n1834, CK => CLK, Q => 
                           n_1211, QN => n14154);
   REGISTERS_reg_16_11_inst : DFF_X1 port map( D => n1833, CK => CLK, Q => 
                           n_1212, QN => n14153);
   REGISTERS_reg_16_10_inst : DFF_X1 port map( D => n1832, CK => CLK, Q => 
                           n_1213, QN => n14152);
   REGISTERS_reg_16_9_inst : DFF_X1 port map( D => n1831, CK => CLK, Q => 
                           n_1214, QN => n14151);
   REGISTERS_reg_16_8_inst : DFF_X1 port map( D => n1830, CK => CLK, Q => 
                           n_1215, QN => n14150);
   REGISTERS_reg_16_7_inst : DFF_X1 port map( D => n1829, CK => CLK, Q => 
                           n_1216, QN => n14149);
   REGISTERS_reg_16_6_inst : DFF_X1 port map( D => n1828, CK => CLK, Q => 
                           n_1217, QN => n14148);
   REGISTERS_reg_16_5_inst : DFF_X1 port map( D => n1827, CK => CLK, Q => 
                           n_1218, QN => n14147);
   REGISTERS_reg_16_4_inst : DFF_X1 port map( D => n1826, CK => CLK, Q => 
                           n_1219, QN => n14146);
   REGISTERS_reg_16_3_inst : DFF_X1 port map( D => n1825, CK => CLK, Q => 
                           n_1220, QN => n14145);
   REGISTERS_reg_16_2_inst : DFF_X1 port map( D => n1824, CK => CLK, Q => 
                           n_1221, QN => n14144);
   REGISTERS_reg_16_1_inst : DFF_X1 port map( D => n1823, CK => CLK, Q => 
                           n_1222, QN => n14143);
   REGISTERS_reg_16_0_inst : DFF_X1 port map( D => n1822, CK => CLK, Q => 
                           n_1223, QN => n14142);
   REGISTERS_reg_17_31_inst : DFF_X1 port map( D => n1821, CK => CLK, Q => 
                           n_1224, QN => n13711);
   REGISTERS_reg_17_30_inst : DFF_X1 port map( D => n1820, CK => CLK, Q => 
                           n_1225, QN => n13710);
   REGISTERS_reg_17_29_inst : DFF_X1 port map( D => n1819, CK => CLK, Q => 
                           n_1226, QN => n13709);
   REGISTERS_reg_17_28_inst : DFF_X1 port map( D => n1818, CK => CLK, Q => 
                           n_1227, QN => n13708);
   REGISTERS_reg_17_27_inst : DFF_X1 port map( D => n1817, CK => CLK, Q => 
                           n_1228, QN => n13707);
   REGISTERS_reg_17_26_inst : DFF_X1 port map( D => n1816, CK => CLK, Q => 
                           n_1229, QN => n13706);
   REGISTERS_reg_17_25_inst : DFF_X1 port map( D => n1815, CK => CLK, Q => 
                           n_1230, QN => n13705);
   REGISTERS_reg_17_24_inst : DFF_X1 port map( D => n1814, CK => CLK, Q => 
                           n_1231, QN => n13704);
   REGISTERS_reg_17_23_inst : DFF_X1 port map( D => n1813, CK => CLK, Q => 
                           n_1232, QN => n13723);
   REGISTERS_reg_17_22_inst : DFF_X1 port map( D => n1812, CK => CLK, Q => 
                           n_1233, QN => n13722);
   REGISTERS_reg_17_21_inst : DFF_X1 port map( D => n1811, CK => CLK, Q => 
                           n_1234, QN => n13721);
   REGISTERS_reg_17_20_inst : DFF_X1 port map( D => n1810, CK => CLK, Q => 
                           n_1235, QN => n13720);
   REGISTERS_reg_17_19_inst : DFF_X1 port map( D => n1809, CK => CLK, Q => 
                           n_1236, QN => n13719);
   REGISTERS_reg_17_18_inst : DFF_X1 port map( D => n1808, CK => CLK, Q => 
                           n_1237, QN => n13718);
   REGISTERS_reg_17_17_inst : DFF_X1 port map( D => n1807, CK => CLK, Q => 
                           n_1238, QN => n13717);
   REGISTERS_reg_17_16_inst : DFF_X1 port map( D => n1806, CK => CLK, Q => 
                           n_1239, QN => n13716);
   REGISTERS_reg_17_15_inst : DFF_X1 port map( D => n1805, CK => CLK, Q => 
                           n_1240, QN => n13715);
   REGISTERS_reg_17_14_inst : DFF_X1 port map( D => n1804, CK => CLK, Q => 
                           n_1241, QN => n13714);
   REGISTERS_reg_17_13_inst : DFF_X1 port map( D => n1803, CK => CLK, Q => 
                           n_1242, QN => n13713);
   REGISTERS_reg_17_12_inst : DFF_X1 port map( D => n1802, CK => CLK, Q => 
                           n_1243, QN => n13712);
   REGISTERS_reg_17_11_inst : DFF_X1 port map( D => n1801, CK => CLK, Q => 
                           n_1244, QN => n13823);
   REGISTERS_reg_17_10_inst : DFF_X1 port map( D => n1800, CK => CLK, Q => 
                           n_1245, QN => n13822);
   REGISTERS_reg_17_9_inst : DFF_X1 port map( D => n1799, CK => CLK, Q => 
                           n_1246, QN => n13821);
   REGISTERS_reg_17_8_inst : DFF_X1 port map( D => n1798, CK => CLK, Q => 
                           n_1247, QN => n13820);
   REGISTERS_reg_17_7_inst : DFF_X1 port map( D => n1797, CK => CLK, Q => 
                           n_1248, QN => n13819);
   REGISTERS_reg_17_6_inst : DFF_X1 port map( D => n1796, CK => CLK, Q => 
                           n_1249, QN => n13818);
   REGISTERS_reg_17_5_inst : DFF_X1 port map( D => n1795, CK => CLK, Q => 
                           n_1250, QN => n13817);
   REGISTERS_reg_17_4_inst : DFF_X1 port map( D => n1794, CK => CLK, Q => 
                           n_1251, QN => n13816);
   REGISTERS_reg_17_3_inst : DFF_X1 port map( D => n1793, CK => CLK, Q => 
                           n_1252, QN => n13815);
   REGISTERS_reg_17_2_inst : DFF_X1 port map( D => n1792, CK => CLK, Q => 
                           n_1253, QN => n13814);
   REGISTERS_reg_17_1_inst : DFF_X1 port map( D => n1791, CK => CLK, Q => 
                           n_1254, QN => n13813);
   REGISTERS_reg_17_0_inst : DFF_X1 port map( D => n1790, CK => CLK, Q => 
                           n_1255, QN => n13812);
   REGISTERS_reg_18_31_inst : DFF_X1 port map( D => n1789, CK => CLK, Q => 
                           n_1256, QN => n13651);
   REGISTERS_reg_18_30_inst : DFF_X1 port map( D => n1788, CK => CLK, Q => 
                           n_1257, QN => n13650);
   REGISTERS_reg_18_29_inst : DFF_X1 port map( D => n1787, CK => CLK, Q => 
                           n_1258, QN => n13649);
   REGISTERS_reg_18_28_inst : DFF_X1 port map( D => n1786, CK => CLK, Q => 
                           n_1259, QN => n13648);
   REGISTERS_reg_18_27_inst : DFF_X1 port map( D => n1785, CK => CLK, Q => 
                           n_1260, QN => n13647);
   REGISTERS_reg_18_26_inst : DFF_X1 port map( D => n1784, CK => CLK, Q => 
                           n_1261, QN => n13646);
   REGISTERS_reg_18_25_inst : DFF_X1 port map( D => n1783, CK => CLK, Q => 
                           n_1262, QN => n13645);
   REGISTERS_reg_18_24_inst : DFF_X1 port map( D => n1782, CK => CLK, Q => 
                           n_1263, QN => n13644);
   REGISTERS_reg_18_23_inst : DFF_X1 port map( D => n1781, CK => CLK, Q => 
                           n_1264, QN => n13671);
   REGISTERS_reg_18_22_inst : DFF_X1 port map( D => n1780, CK => CLK, Q => 
                           n_1265, QN => n13670);
   REGISTERS_reg_18_21_inst : DFF_X1 port map( D => n1779, CK => CLK, Q => 
                           n_1266, QN => n13669);
   REGISTERS_reg_18_20_inst : DFF_X1 port map( D => n1778, CK => CLK, Q => 
                           n_1267, QN => n13668);
   REGISTERS_reg_18_19_inst : DFF_X1 port map( D => n1777, CK => CLK, Q => 
                           n_1268, QN => n13667);
   REGISTERS_reg_18_18_inst : DFF_X1 port map( D => n1776, CK => CLK, Q => 
                           n_1269, QN => n13666);
   REGISTERS_reg_18_17_inst : DFF_X1 port map( D => n1775, CK => CLK, Q => 
                           n_1270, QN => n13665);
   REGISTERS_reg_18_16_inst : DFF_X1 port map( D => n1774, CK => CLK, Q => 
                           n_1271, QN => n13664);
   REGISTERS_reg_18_15_inst : DFF_X1 port map( D => n1773, CK => CLK, Q => 
                           n_1272, QN => n13663);
   REGISTERS_reg_18_14_inst : DFF_X1 port map( D => n1772, CK => CLK, Q => 
                           n_1273, QN => n13662);
   REGISTERS_reg_18_13_inst : DFF_X1 port map( D => n1771, CK => CLK, Q => 
                           n_1274, QN => n13661);
   REGISTERS_reg_18_12_inst : DFF_X1 port map( D => n1770, CK => CLK, Q => 
                           n_1275, QN => n13660);
   REGISTERS_reg_18_11_inst : DFF_X1 port map( D => n1769, CK => CLK, Q => 
                           n_1276, QN => n13739);
   REGISTERS_reg_18_10_inst : DFF_X1 port map( D => n1768, CK => CLK, Q => 
                           n_1277, QN => n13738);
   REGISTERS_reg_18_9_inst : DFF_X1 port map( D => n1767, CK => CLK, Q => 
                           n_1278, QN => n13737);
   REGISTERS_reg_18_8_inst : DFF_X1 port map( D => n1766, CK => CLK, Q => 
                           n_1279, QN => n13736);
   REGISTERS_reg_18_7_inst : DFF_X1 port map( D => n1765, CK => CLK, Q => 
                           n_1280, QN => n13735);
   REGISTERS_reg_18_6_inst : DFF_X1 port map( D => n1764, CK => CLK, Q => 
                           n_1281, QN => n13734);
   REGISTERS_reg_18_5_inst : DFF_X1 port map( D => n1763, CK => CLK, Q => 
                           n_1282, QN => n13733);
   REGISTERS_reg_18_4_inst : DFF_X1 port map( D => n1762, CK => CLK, Q => 
                           n_1283, QN => n13732);
   REGISTERS_reg_18_3_inst : DFF_X1 port map( D => n1761, CK => CLK, Q => 
                           n_1284, QN => n13731);
   REGISTERS_reg_18_2_inst : DFF_X1 port map( D => n1760, CK => CLK, Q => 
                           n_1285, QN => n13730);
   REGISTERS_reg_18_1_inst : DFF_X1 port map( D => n1759, CK => CLK, Q => 
                           n_1286, QN => n13729);
   REGISTERS_reg_18_0_inst : DFF_X1 port map( D => n1758, CK => CLK, Q => 
                           n_1287, QN => n13728);
   REGISTERS_reg_19_31_inst : DFF_X1 port map( D => n1757, CK => CLK, Q => 
                           n_1288, QN => n13907);
   REGISTERS_reg_19_30_inst : DFF_X1 port map( D => n1756, CK => CLK, Q => 
                           n_1289, QN => n13905);
   REGISTERS_reg_19_29_inst : DFF_X1 port map( D => n1755, CK => CLK, Q => 
                           n_1290, QN => n13903);
   REGISTERS_reg_19_28_inst : DFF_X1 port map( D => n1754, CK => CLK, Q => 
                           n_1291, QN => n13901);
   REGISTERS_reg_19_27_inst : DFF_X1 port map( D => n1753, CK => CLK, Q => 
                           n_1292, QN => n13899);
   REGISTERS_reg_19_26_inst : DFF_X1 port map( D => n1752, CK => CLK, Q => 
                           n_1293, QN => n13897);
   REGISTERS_reg_19_25_inst : DFF_X1 port map( D => n1751, CK => CLK, Q => 
                           n_1294, QN => n13895);
   REGISTERS_reg_19_24_inst : DFF_X1 port map( D => n1750, CK => CLK, Q => 
                           n_1295, QN => n13893);
   REGISTERS_reg_19_23_inst : DFF_X1 port map( D => n1749, CK => CLK, Q => 
                           n_1296, QN => n14193);
   REGISTERS_reg_19_22_inst : DFF_X1 port map( D => n1748, CK => CLK, Q => 
                           n_1297, QN => n14191);
   REGISTERS_reg_19_21_inst : DFF_X1 port map( D => n1747, CK => CLK, Q => 
                           n_1298, QN => n14189);
   REGISTERS_reg_19_20_inst : DFF_X1 port map( D => n1746, CK => CLK, Q => 
                           n_1299, QN => n14187);
   REGISTERS_reg_19_19_inst : DFF_X1 port map( D => n1745, CK => CLK, Q => 
                           n_1300, QN => n14185);
   REGISTERS_reg_19_18_inst : DFF_X1 port map( D => n1744, CK => CLK, Q => 
                           n_1301, QN => n14183);
   REGISTERS_reg_19_17_inst : DFF_X1 port map( D => n1743, CK => CLK, Q => 
                           n_1302, QN => n14181);
   REGISTERS_reg_19_16_inst : DFF_X1 port map( D => n1742, CK => CLK, Q => 
                           n_1303, QN => n14179);
   REGISTERS_reg_19_15_inst : DFF_X1 port map( D => n1741, CK => CLK, Q => 
                           n_1304, QN => n14177);
   REGISTERS_reg_19_14_inst : DFF_X1 port map( D => n1740, CK => CLK, Q => 
                           n_1305, QN => n14175);
   REGISTERS_reg_19_13_inst : DFF_X1 port map( D => n1739, CK => CLK, Q => 
                           n_1306, QN => n14173);
   REGISTERS_reg_19_12_inst : DFF_X1 port map( D => n1738, CK => CLK, Q => 
                           n_1307, QN => n14171);
   REGISTERS_reg_19_11_inst : DFF_X1 port map( D => n1737, CK => CLK, Q => 
                           n_1308, QN => n14169);
   REGISTERS_reg_19_10_inst : DFF_X1 port map( D => n1736, CK => CLK, Q => 
                           n_1309, QN => n14168);
   REGISTERS_reg_19_9_inst : DFF_X1 port map( D => n1735, CK => CLK, Q => 
                           n_1310, QN => n14167);
   REGISTERS_reg_19_8_inst : DFF_X1 port map( D => n1734, CK => CLK, Q => 
                           n_1311, QN => n14166);
   REGISTERS_reg_19_7_inst : DFF_X1 port map( D => n1733, CK => CLK, Q => 
                           n_1312, QN => n14225);
   REGISTERS_reg_19_6_inst : DFF_X1 port map( D => n1732, CK => CLK, Q => 
                           n_1313, QN => n14224);
   REGISTERS_reg_19_5_inst : DFF_X1 port map( D => n1731, CK => CLK, Q => 
                           n_1314, QN => n14223);
   REGISTERS_reg_19_4_inst : DFF_X1 port map( D => n1730, CK => CLK, Q => 
                           n_1315, QN => n14222);
   REGISTERS_reg_19_3_inst : DFF_X1 port map( D => n1729, CK => CLK, Q => 
                           n_1316, QN => n14221);
   REGISTERS_reg_19_2_inst : DFF_X1 port map( D => n1728, CK => CLK, Q => 
                           n_1317, QN => n14220);
   REGISTERS_reg_19_1_inst : DFF_X1 port map( D => n1727, CK => CLK, Q => 
                           n_1318, QN => n14219);
   REGISTERS_reg_19_0_inst : DFF_X1 port map( D => n1726, CK => CLK, Q => 
                           n_1319, QN => n14218);
   REGISTERS_reg_20_31_inst : DFF_X1 port map( D => n1725, CK => CLK, Q => 
                           n_1320, QN => n13811);
   REGISTERS_reg_20_30_inst : DFF_X1 port map( D => n1724, CK => CLK, Q => 
                           n_1321, QN => n13810);
   REGISTERS_reg_20_29_inst : DFF_X1 port map( D => n1723, CK => CLK, Q => 
                           n_1322, QN => n13809);
   REGISTERS_reg_20_28_inst : DFF_X1 port map( D => n1722, CK => CLK, Q => 
                           n_1323, QN => n13808);
   REGISTERS_reg_20_27_inst : DFF_X1 port map( D => n1721, CK => CLK, Q => 
                           n_1324, QN => n13807);
   REGISTERS_reg_20_26_inst : DFF_X1 port map( D => n1720, CK => CLK, Q => 
                           n_1325, QN => n13806);
   REGISTERS_reg_20_25_inst : DFF_X1 port map( D => n1719, CK => CLK, Q => 
                           n_1326, QN => n13805);
   REGISTERS_reg_20_24_inst : DFF_X1 port map( D => n1718, CK => CLK, Q => 
                           n_1327, QN => n13804);
   REGISTERS_reg_20_23_inst : DFF_X1 port map( D => n1717, CK => CLK, Q => 
                           n_1328, QN => n14069);
   REGISTERS_reg_20_22_inst : DFF_X1 port map( D => n1716, CK => CLK, Q => 
                           n_1329, QN => n14068);
   REGISTERS_reg_20_21_inst : DFF_X1 port map( D => n1715, CK => CLK, Q => 
                           n_1330, QN => n14067);
   REGISTERS_reg_20_20_inst : DFF_X1 port map( D => n1714, CK => CLK, Q => 
                           n_1331, QN => n14066);
   REGISTERS_reg_20_19_inst : DFF_X1 port map( D => n1713, CK => CLK, Q => 
                           n_1332, QN => n14065);
   REGISTERS_reg_20_18_inst : DFF_X1 port map( D => n1712, CK => CLK, Q => 
                           n_1333, QN => n14064);
   REGISTERS_reg_20_17_inst : DFF_X1 port map( D => n1711, CK => CLK, Q => 
                           n_1334, QN => n14063);
   REGISTERS_reg_20_16_inst : DFF_X1 port map( D => n1710, CK => CLK, Q => 
                           n_1335, QN => n14062);
   REGISTERS_reg_20_15_inst : DFF_X1 port map( D => n1709, CK => CLK, Q => 
                           n_1336, QN => n14061);
   REGISTERS_reg_20_14_inst : DFF_X1 port map( D => n1708, CK => CLK, Q => 
                           n_1337, QN => n14060);
   REGISTERS_reg_20_13_inst : DFF_X1 port map( D => n1707, CK => CLK, Q => 
                           n_1338, QN => n14059);
   REGISTERS_reg_20_12_inst : DFF_X1 port map( D => n1706, CK => CLK, Q => 
                           n_1339, QN => n14058);
   REGISTERS_reg_20_11_inst : DFF_X1 port map( D => n1705, CK => CLK, Q => 
                           n_1340, QN => n14057);
   REGISTERS_reg_20_10_inst : DFF_X1 port map( D => n1704, CK => CLK, Q => 
                           n_1341, QN => n14056);
   REGISTERS_reg_20_9_inst : DFF_X1 port map( D => n1703, CK => CLK, Q => 
                           n_1342, QN => n14055);
   REGISTERS_reg_20_8_inst : DFF_X1 port map( D => n1702, CK => CLK, Q => 
                           n_1343, QN => n14054);
   REGISTERS_reg_20_7_inst : DFF_X1 port map( D => n1701, CK => CLK, Q => 
                           n_1344, QN => n14053);
   REGISTERS_reg_20_6_inst : DFF_X1 port map( D => n1700, CK => CLK, Q => 
                           n_1345, QN => n14052);
   REGISTERS_reg_20_5_inst : DFF_X1 port map( D => n1699, CK => CLK, Q => 
                           n_1346, QN => n14051);
   REGISTERS_reg_20_4_inst : DFF_X1 port map( D => n1698, CK => CLK, Q => 
                           n_1347, QN => n14050);
   REGISTERS_reg_20_3_inst : DFF_X1 port map( D => n1697, CK => CLK, Q => 
                           n_1348, QN => n14049);
   REGISTERS_reg_20_2_inst : DFF_X1 port map( D => n1696, CK => CLK, Q => 
                           n_1349, QN => n14048);
   REGISTERS_reg_20_1_inst : DFF_X1 port map( D => n1695, CK => CLK, Q => 
                           n_1350, QN => n14047);
   REGISTERS_reg_20_0_inst : DFF_X1 port map( D => n1694, CK => CLK, Q => 
                           n_1351, QN => n14046);
   REGISTERS_reg_21_31_inst : DFF_X1 port map( D => n1693, CK => CLK, Q => 
                           n_1352, QN => n13891);
   REGISTERS_reg_21_30_inst : DFF_X1 port map( D => n1692, CK => CLK, Q => 
                           n_1353, QN => n13890);
   REGISTERS_reg_21_29_inst : DFF_X1 port map( D => n1691, CK => CLK, Q => 
                           n_1354, QN => n13889);
   REGISTERS_reg_21_28_inst : DFF_X1 port map( D => n1690, CK => CLK, Q => 
                           n_1355, QN => n13888);
   REGISTERS_reg_21_27_inst : DFF_X1 port map( D => n1689, CK => CLK, Q => 
                           n_1356, QN => n13887);
   REGISTERS_reg_21_26_inst : DFF_X1 port map( D => n1688, CK => CLK, Q => 
                           n_1357, QN => n13886);
   REGISTERS_reg_21_25_inst : DFF_X1 port map( D => n1687, CK => CLK, Q => 
                           n_1358, QN => n13885);
   REGISTERS_reg_21_24_inst : DFF_X1 port map( D => n1686, CK => CLK, Q => 
                           n_1359, QN => n13884);
   REGISTERS_reg_21_23_inst : DFF_X1 port map( D => n1685, CK => CLK, Q => 
                           n_1360, QN => n14217);
   REGISTERS_reg_21_22_inst : DFF_X1 port map( D => n1684, CK => CLK, Q => 
                           n_1361, QN => n14216);
   REGISTERS_reg_21_21_inst : DFF_X1 port map( D => n1683, CK => CLK, Q => 
                           n_1362, QN => n14215);
   REGISTERS_reg_21_20_inst : DFF_X1 port map( D => n1682, CK => CLK, Q => 
                           n_1363, QN => n14214);
   REGISTERS_reg_21_19_inst : DFF_X1 port map( D => n1681, CK => CLK, Q => 
                           n_1364, QN => n14213);
   REGISTERS_reg_21_18_inst : DFF_X1 port map( D => n1680, CK => CLK, Q => 
                           n_1365, QN => n14212);
   REGISTERS_reg_21_17_inst : DFF_X1 port map( D => n1679, CK => CLK, Q => 
                           n_1366, QN => n14211);
   REGISTERS_reg_21_16_inst : DFF_X1 port map( D => n1678, CK => CLK, Q => 
                           n_1367, QN => n14210);
   REGISTERS_reg_21_15_inst : DFF_X1 port map( D => n1677, CK => CLK, Q => 
                           n_1368, QN => n14209);
   REGISTERS_reg_21_14_inst : DFF_X1 port map( D => n1676, CK => CLK, Q => 
                           n_1369, QN => n14208);
   REGISTERS_reg_21_13_inst : DFF_X1 port map( D => n1675, CK => CLK, Q => 
                           n_1370, QN => n14207);
   REGISTERS_reg_21_12_inst : DFF_X1 port map( D => n1674, CK => CLK, Q => 
                           n_1371, QN => n14206);
   REGISTERS_reg_21_11_inst : DFF_X1 port map( D => n1673, CK => CLK, Q => 
                           n_1372, QN => n14205);
   REGISTERS_reg_21_10_inst : DFF_X1 port map( D => n1672, CK => CLK, Q => 
                           n_1373, QN => n14204);
   REGISTERS_reg_21_9_inst : DFF_X1 port map( D => n1671, CK => CLK, Q => 
                           n_1374, QN => n14203);
   REGISTERS_reg_21_8_inst : DFF_X1 port map( D => n1670, CK => CLK, Q => 
                           n_1375, QN => n14202);
   REGISTERS_reg_21_7_inst : DFF_X1 port map( D => n1669, CK => CLK, Q => 
                           n_1376, QN => n14201);
   REGISTERS_reg_21_6_inst : DFF_X1 port map( D => n1668, CK => CLK, Q => 
                           n_1377, QN => n14200);
   REGISTERS_reg_21_5_inst : DFF_X1 port map( D => n1667, CK => CLK, Q => 
                           n_1378, QN => n14199);
   REGISTERS_reg_21_4_inst : DFF_X1 port map( D => n1666, CK => CLK, Q => 
                           n_1379, QN => n14198);
   REGISTERS_reg_21_3_inst : DFF_X1 port map( D => n1665, CK => CLK, Q => 
                           n_1380, QN => n14197);
   REGISTERS_reg_21_2_inst : DFF_X1 port map( D => n1664, CK => CLK, Q => 
                           n_1381, QN => n14196);
   REGISTERS_reg_21_1_inst : DFF_X1 port map( D => n1663, CK => CLK, Q => 
                           n_1382, QN => n14195);
   REGISTERS_reg_21_0_inst : DFF_X1 port map( D => n1662, CK => CLK, Q => 
                           n_1383, QN => n14194);
   REGISTERS_reg_22_31_inst : DFF_X1 port map( D => n1661, CK => CLK, Q => 
                           n_1384, QN => n13691);
   REGISTERS_reg_22_30_inst : DFF_X1 port map( D => n1660, CK => CLK, Q => 
                           n_1385, QN => n13690);
   REGISTERS_reg_22_29_inst : DFF_X1 port map( D => n1659, CK => CLK, Q => 
                           n_1386, QN => n13689);
   REGISTERS_reg_22_28_inst : DFF_X1 port map( D => n1658, CK => CLK, Q => 
                           n_1387, QN => n13688);
   REGISTERS_reg_22_27_inst : DFF_X1 port map( D => n1657, CK => CLK, Q => 
                           n_1388, QN => n13687);
   REGISTERS_reg_22_26_inst : DFF_X1 port map( D => n1656, CK => CLK, Q => 
                           n_1389, QN => n13686);
   REGISTERS_reg_22_25_inst : DFF_X1 port map( D => n1655, CK => CLK, Q => 
                           n_1390, QN => n13685);
   REGISTERS_reg_22_24_inst : DFF_X1 port map( D => n1654, CK => CLK, Q => 
                           n_1391, QN => n13684);
   REGISTERS_reg_22_23_inst : DFF_X1 port map( D => n1653, CK => CLK, Q => 
                           n_1392, QN => n13703);
   REGISTERS_reg_22_22_inst : DFF_X1 port map( D => n1652, CK => CLK, Q => 
                           n_1393, QN => n13702);
   REGISTERS_reg_22_21_inst : DFF_X1 port map( D => n1651, CK => CLK, Q => 
                           n_1394, QN => n13701);
   REGISTERS_reg_22_20_inst : DFF_X1 port map( D => n1650, CK => CLK, Q => 
                           n_1395, QN => n13700);
   REGISTERS_reg_22_19_inst : DFF_X1 port map( D => n1649, CK => CLK, Q => 
                           n_1396, QN => n13699);
   REGISTERS_reg_22_18_inst : DFF_X1 port map( D => n1648, CK => CLK, Q => 
                           n_1397, QN => n13698);
   REGISTERS_reg_22_17_inst : DFF_X1 port map( D => n1647, CK => CLK, Q => 
                           n_1398, QN => n13697);
   REGISTERS_reg_22_16_inst : DFF_X1 port map( D => n1646, CK => CLK, Q => 
                           n_1399, QN => n13696);
   REGISTERS_reg_22_15_inst : DFF_X1 port map( D => n1645, CK => CLK, Q => 
                           n_1400, QN => n13695);
   REGISTERS_reg_22_14_inst : DFF_X1 port map( D => n1644, CK => CLK, Q => 
                           n_1401, QN => n13694);
   REGISTERS_reg_22_13_inst : DFF_X1 port map( D => n1643, CK => CLK, Q => 
                           n_1402, QN => n13693);
   REGISTERS_reg_22_12_inst : DFF_X1 port map( D => n1642, CK => CLK, Q => 
                           n_1403, QN => n13692);
   REGISTERS_reg_22_11_inst : DFF_X1 port map( D => n1641, CK => CLK, Q => 
                           n_1404, QN => n13803);
   REGISTERS_reg_22_10_inst : DFF_X1 port map( D => n1640, CK => CLK, Q => 
                           n_1405, QN => n13802);
   REGISTERS_reg_22_9_inst : DFF_X1 port map( D => n1639, CK => CLK, Q => 
                           n_1406, QN => n13801);
   REGISTERS_reg_22_8_inst : DFF_X1 port map( D => n1638, CK => CLK, Q => 
                           n_1407, QN => n13800);
   REGISTERS_reg_22_7_inst : DFF_X1 port map( D => n1637, CK => CLK, Q => 
                           n_1408, QN => n13799);
   REGISTERS_reg_22_6_inst : DFF_X1 port map( D => n1636, CK => CLK, Q => 
                           n_1409, QN => n13798);
   REGISTERS_reg_22_5_inst : DFF_X1 port map( D => n1635, CK => CLK, Q => 
                           n_1410, QN => n13797);
   REGISTERS_reg_22_4_inst : DFF_X1 port map( D => n1634, CK => CLK, Q => 
                           n_1411, QN => n13796);
   REGISTERS_reg_22_3_inst : DFF_X1 port map( D => n1633, CK => CLK, Q => 
                           n_1412, QN => n13795);
   REGISTERS_reg_22_2_inst : DFF_X1 port map( D => n1632, CK => CLK, Q => 
                           n_1413, QN => n13794);
   REGISTERS_reg_22_1_inst : DFF_X1 port map( D => n1631, CK => CLK, Q => 
                           n_1414, QN => n13793);
   REGISTERS_reg_22_0_inst : DFF_X1 port map( D => n1630, CK => CLK, Q => 
                           n_1415, QN => n13792);
   REGISTERS_reg_23_31_inst : DFF_X1 port map( D => n1629, CK => CLK, Q => 
                           n_1416, QN => n13906);
   REGISTERS_reg_23_30_inst : DFF_X1 port map( D => n1628, CK => CLK, Q => 
                           n_1417, QN => n13904);
   REGISTERS_reg_23_29_inst : DFF_X1 port map( D => n1627, CK => CLK, Q => 
                           n_1418, QN => n13902);
   REGISTERS_reg_23_28_inst : DFF_X1 port map( D => n1626, CK => CLK, Q => 
                           n_1419, QN => n13900);
   REGISTERS_reg_23_27_inst : DFF_X1 port map( D => n1625, CK => CLK, Q => 
                           n_1420, QN => n13898);
   REGISTERS_reg_23_26_inst : DFF_X1 port map( D => n1624, CK => CLK, Q => 
                           n_1421, QN => n13896);
   REGISTERS_reg_23_25_inst : DFF_X1 port map( D => n1623, CK => CLK, Q => 
                           n_1422, QN => n13894);
   REGISTERS_reg_23_24_inst : DFF_X1 port map( D => n1622, CK => CLK, Q => 
                           n_1423, QN => n13892);
   REGISTERS_reg_23_23_inst : DFF_X1 port map( D => n1621, CK => CLK, Q => 
                           n_1424, QN => n14192);
   REGISTERS_reg_23_22_inst : DFF_X1 port map( D => n1620, CK => CLK, Q => 
                           n_1425, QN => n14190);
   REGISTERS_reg_23_21_inst : DFF_X1 port map( D => n1619, CK => CLK, Q => 
                           n_1426, QN => n14188);
   REGISTERS_reg_23_20_inst : DFF_X1 port map( D => n1618, CK => CLK, Q => 
                           n_1427, QN => n14186);
   REGISTERS_reg_23_19_inst : DFF_X1 port map( D => n1617, CK => CLK, Q => 
                           n_1428, QN => n14184);
   REGISTERS_reg_23_18_inst : DFF_X1 port map( D => n1616, CK => CLK, Q => 
                           n_1429, QN => n14182);
   REGISTERS_reg_23_17_inst : DFF_X1 port map( D => n1615, CK => CLK, Q => 
                           n_1430, QN => n14180);
   REGISTERS_reg_23_16_inst : DFF_X1 port map( D => n1614, CK => CLK, Q => 
                           n_1431, QN => n14178);
   REGISTERS_reg_23_15_inst : DFF_X1 port map( D => n1613, CK => CLK, Q => 
                           n_1432, QN => n14176);
   REGISTERS_reg_23_14_inst : DFF_X1 port map( D => n1612, CK => CLK, Q => 
                           n_1433, QN => n14174);
   REGISTERS_reg_23_13_inst : DFF_X1 port map( D => n1611, CK => CLK, Q => 
                           n_1434, QN => n14172);
   REGISTERS_reg_23_12_inst : DFF_X1 port map( D => n1610, CK => CLK, Q => 
                           n_1435, QN => n14170);
   REGISTERS_reg_23_11_inst : DFF_X1 port map( D => n1609, CK => CLK, Q => 
                           n_1436, QN => n13883);
   REGISTERS_reg_23_10_inst : DFF_X1 port map( D => n1608, CK => CLK, Q => 
                           n_1437, QN => n13882);
   REGISTERS_reg_23_9_inst : DFF_X1 port map( D => n1607, CK => CLK, Q => 
                           n_1438, QN => n13881);
   REGISTERS_reg_23_8_inst : DFF_X1 port map( D => n1606, CK => CLK, Q => 
                           n_1439, QN => n13880);
   REGISTERS_reg_23_7_inst : DFF_X1 port map( D => n1605, CK => CLK, Q => 
                           n_1440, QN => n13915);
   REGISTERS_reg_23_6_inst : DFF_X1 port map( D => n1604, CK => CLK, Q => 
                           n_1441, QN => n13914);
   REGISTERS_reg_23_5_inst : DFF_X1 port map( D => n1603, CK => CLK, Q => 
                           n_1442, QN => n13913);
   REGISTERS_reg_23_4_inst : DFF_X1 port map( D => n1602, CK => CLK, Q => 
                           n_1443, QN => n13912);
   REGISTERS_reg_23_3_inst : DFF_X1 port map( D => n1601, CK => CLK, Q => 
                           n_1444, QN => n13911);
   REGISTERS_reg_23_2_inst : DFF_X1 port map( D => n1600, CK => CLK, Q => 
                           n_1445, QN => n13910);
   REGISTERS_reg_23_1_inst : DFF_X1 port map( D => n1599, CK => CLK, Q => 
                           n_1446, QN => n13909);
   REGISTERS_reg_23_0_inst : DFF_X1 port map( D => n1598, CK => CLK, Q => 
                           n_1447, QN => n13908);
   REGISTERS_reg_24_31_inst : DFF_X1 port map( D => n1597, CK => CLK, Q => 
                           n13947, QN => n9404);
   REGISTERS_reg_24_30_inst : DFF_X1 port map( D => n1596, CK => CLK, Q => 
                           n13946, QN => n9405);
   REGISTERS_reg_24_29_inst : DFF_X1 port map( D => n1595, CK => CLK, Q => 
                           n13945, QN => n9406);
   REGISTERS_reg_24_28_inst : DFF_X1 port map( D => n1594, CK => CLK, Q => 
                           n13944, QN => n9407);
   REGISTERS_reg_24_27_inst : DFF_X1 port map( D => n1593, CK => CLK, Q => 
                           n13943, QN => n9408);
   REGISTERS_reg_24_26_inst : DFF_X1 port map( D => n1592, CK => CLK, Q => 
                           n13942, QN => n9409);
   REGISTERS_reg_24_25_inst : DFF_X1 port map( D => n1591, CK => CLK, Q => 
                           n13941, QN => n9410);
   REGISTERS_reg_24_24_inst : DFF_X1 port map( D => n1590, CK => CLK, Q => 
                           n13940, QN => n9411);
   REGISTERS_reg_24_23_inst : DFF_X1 port map( D => n1589, CK => CLK, Q => 
                           n13939, QN => n9412);
   REGISTERS_reg_24_22_inst : DFF_X1 port map( D => n1588, CK => CLK, Q => 
                           n13938, QN => n9413);
   REGISTERS_reg_24_21_inst : DFF_X1 port map( D => n1587, CK => CLK, Q => 
                           n13937, QN => n9414);
   REGISTERS_reg_24_20_inst : DFF_X1 port map( D => n1586, CK => CLK, Q => 
                           n13936, QN => n9415);
   REGISTERS_reg_24_19_inst : DFF_X1 port map( D => n1585, CK => CLK, Q => 
                           n13935, QN => n9416);
   REGISTERS_reg_24_18_inst : DFF_X1 port map( D => n1584, CK => CLK, Q => 
                           n13934, QN => n9417);
   REGISTERS_reg_24_17_inst : DFF_X1 port map( D => n1583, CK => CLK, Q => 
                           n13933, QN => n9418);
   REGISTERS_reg_24_16_inst : DFF_X1 port map( D => n1582, CK => CLK, Q => 
                           n13932, QN => n9419);
   REGISTERS_reg_24_15_inst : DFF_X1 port map( D => n1581, CK => CLK, Q => 
                           n13931, QN => n9420);
   REGISTERS_reg_24_14_inst : DFF_X1 port map( D => n1580, CK => CLK, Q => 
                           n13930, QN => n9421);
   REGISTERS_reg_24_13_inst : DFF_X1 port map( D => n1579, CK => CLK, Q => 
                           n13929, QN => n9422);
   REGISTERS_reg_24_12_inst : DFF_X1 port map( D => n1578, CK => CLK, Q => 
                           n13928, QN => n9423);
   REGISTERS_reg_24_11_inst : DFF_X1 port map( D => n1577, CK => CLK, Q => 
                           n13927, QN => n9424);
   REGISTERS_reg_24_10_inst : DFF_X1 port map( D => n1576, CK => CLK, Q => 
                           n13926, QN => n9425);
   REGISTERS_reg_24_9_inst : DFF_X1 port map( D => n1575, CK => CLK, Q => 
                           n13925, QN => n9426);
   REGISTERS_reg_24_8_inst : DFF_X1 port map( D => n1574, CK => CLK, Q => 
                           n13924, QN => n9427);
   REGISTERS_reg_24_7_inst : DFF_X1 port map( D => n1573, CK => CLK, Q => 
                           n13923, QN => n9428);
   REGISTERS_reg_24_6_inst : DFF_X1 port map( D => n1572, CK => CLK, Q => 
                           n13922, QN => n9429);
   REGISTERS_reg_24_5_inst : DFF_X1 port map( D => n1571, CK => CLK, Q => 
                           n13921, QN => n9430);
   REGISTERS_reg_24_4_inst : DFF_X1 port map( D => n1570, CK => CLK, Q => 
                           n13920, QN => n9431);
   REGISTERS_reg_24_3_inst : DFF_X1 port map( D => n1569, CK => CLK, Q => 
                           n13919, QN => n9432);
   REGISTERS_reg_24_2_inst : DFF_X1 port map( D => n1568, CK => CLK, Q => 
                           n13918, QN => n9433);
   REGISTERS_reg_24_1_inst : DFF_X1 port map( D => n1567, CK => CLK, Q => 
                           n13917, QN => n9434);
   REGISTERS_reg_24_0_inst : DFF_X1 port map( D => n1566, CK => CLK, Q => 
                           n13916, QN => n9435);
   REGISTERS_reg_25_31_inst : DFF_X1 port map( D => n1565, CK => CLK, Q => 
                           n14257, QN => n9436);
   REGISTERS_reg_25_30_inst : DFF_X1 port map( D => n1564, CK => CLK, Q => 
                           n14256, QN => n9437);
   REGISTERS_reg_25_29_inst : DFF_X1 port map( D => n1563, CK => CLK, Q => 
                           n14255, QN => n9438);
   REGISTERS_reg_25_28_inst : DFF_X1 port map( D => n1562, CK => CLK, Q => 
                           n14254, QN => n9439);
   REGISTERS_reg_25_27_inst : DFF_X1 port map( D => n1561, CK => CLK, Q => 
                           n14253, QN => n9440);
   REGISTERS_reg_25_26_inst : DFF_X1 port map( D => n1560, CK => CLK, Q => 
                           n14252, QN => n9441);
   REGISTERS_reg_25_25_inst : DFF_X1 port map( D => n1559, CK => CLK, Q => 
                           n14251, QN => n9442);
   REGISTERS_reg_25_24_inst : DFF_X1 port map( D => n1558, CK => CLK, Q => 
                           n14250, QN => n9443);
   REGISTERS_reg_25_23_inst : DFF_X1 port map( D => n1557, CK => CLK, Q => 
                           n14249, QN => n9444);
   REGISTERS_reg_25_22_inst : DFF_X1 port map( D => n1556, CK => CLK, Q => 
                           n14248, QN => n9445);
   REGISTERS_reg_25_21_inst : DFF_X1 port map( D => n1555, CK => CLK, Q => 
                           n14247, QN => n9446);
   REGISTERS_reg_25_20_inst : DFF_X1 port map( D => n1554, CK => CLK, Q => 
                           n14246, QN => n9447);
   REGISTERS_reg_25_19_inst : DFF_X1 port map( D => n1553, CK => CLK, Q => 
                           n14245, QN => n9448);
   REGISTERS_reg_25_18_inst : DFF_X1 port map( D => n1552, CK => CLK, Q => 
                           n14244, QN => n9449);
   REGISTERS_reg_25_17_inst : DFF_X1 port map( D => n1551, CK => CLK, Q => 
                           n14243, QN => n9450);
   REGISTERS_reg_25_16_inst : DFF_X1 port map( D => n1550, CK => CLK, Q => 
                           n14242, QN => n9451);
   REGISTERS_reg_25_15_inst : DFF_X1 port map( D => n1549, CK => CLK, Q => 
                           n14241, QN => n9452);
   REGISTERS_reg_25_14_inst : DFF_X1 port map( D => n1548, CK => CLK, Q => 
                           n14240, QN => n9453);
   REGISTERS_reg_25_13_inst : DFF_X1 port map( D => n1547, CK => CLK, Q => 
                           n14239, QN => n9454);
   REGISTERS_reg_25_12_inst : DFF_X1 port map( D => n1546, CK => CLK, Q => 
                           n14238, QN => n9455);
   REGISTERS_reg_25_11_inst : DFF_X1 port map( D => n1545, CK => CLK, Q => 
                           n14237, QN => n9456);
   REGISTERS_reg_25_10_inst : DFF_X1 port map( D => n1544, CK => CLK, Q => 
                           n14236, QN => n9457);
   REGISTERS_reg_25_9_inst : DFF_X1 port map( D => n1543, CK => CLK, Q => 
                           n14235, QN => n9458);
   REGISTERS_reg_25_8_inst : DFF_X1 port map( D => n1542, CK => CLK, Q => 
                           n14234, QN => n9459);
   REGISTERS_reg_25_7_inst : DFF_X1 port map( D => n1541, CK => CLK, Q => 
                           n14233, QN => n9460);
   REGISTERS_reg_25_6_inst : DFF_X1 port map( D => n1540, CK => CLK, Q => 
                           n14232, QN => n9461);
   REGISTERS_reg_25_5_inst : DFF_X1 port map( D => n1539, CK => CLK, Q => 
                           n14231, QN => n9462);
   REGISTERS_reg_25_4_inst : DFF_X1 port map( D => n1538, CK => CLK, Q => 
                           n14230, QN => n9463);
   REGISTERS_reg_25_3_inst : DFF_X1 port map( D => n1537, CK => CLK, Q => 
                           n14229, QN => n9464);
   REGISTERS_reg_25_2_inst : DFF_X1 port map( D => n1536, CK => CLK, Q => 
                           n14228, QN => n9465);
   REGISTERS_reg_25_1_inst : DFF_X1 port map( D => n1535, CK => CLK, Q => 
                           n14227, QN => n9466);
   REGISTERS_reg_25_0_inst : DFF_X1 port map( D => n1534, CK => CLK, Q => 
                           n14226, QN => n9467);
   REGISTERS_reg_26_31_inst : DFF_X1 port map( D => n1533, CK => CLK, Q => 
                           n14353, QN => n9468);
   REGISTERS_reg_26_30_inst : DFF_X1 port map( D => n1532, CK => CLK, Q => 
                           n14352, QN => n9469);
   REGISTERS_reg_26_29_inst : DFF_X1 port map( D => n1531, CK => CLK, Q => 
                           n14351, QN => n9470);
   REGISTERS_reg_26_28_inst : DFF_X1 port map( D => n1530, CK => CLK, Q => 
                           n14350, QN => n9471);
   REGISTERS_reg_26_27_inst : DFF_X1 port map( D => n1529, CK => CLK, Q => 
                           n14349, QN => n9472);
   REGISTERS_reg_26_26_inst : DFF_X1 port map( D => n1528, CK => CLK, Q => 
                           n14348, QN => n9473);
   REGISTERS_reg_26_25_inst : DFF_X1 port map( D => n1527, CK => CLK, Q => 
                           n14347, QN => n9474);
   REGISTERS_reg_26_24_inst : DFF_X1 port map( D => n1526, CK => CLK, Q => 
                           n14346, QN => n9475);
   REGISTERS_reg_26_23_inst : DFF_X1 port map( D => n1525, CK => CLK, Q => 
                           n14345, QN => n9476);
   REGISTERS_reg_26_22_inst : DFF_X1 port map( D => n1524, CK => CLK, Q => 
                           n14344, QN => n9477);
   REGISTERS_reg_26_21_inst : DFF_X1 port map( D => n1523, CK => CLK, Q => 
                           n14343, QN => n9478);
   REGISTERS_reg_26_20_inst : DFF_X1 port map( D => n1522, CK => CLK, Q => 
                           n14342, QN => n9479);
   REGISTERS_reg_26_19_inst : DFF_X1 port map( D => n1521, CK => CLK, Q => 
                           n14341, QN => n9480);
   REGISTERS_reg_26_18_inst : DFF_X1 port map( D => n1520, CK => CLK, Q => 
                           n14340, QN => n9481);
   REGISTERS_reg_26_17_inst : DFF_X1 port map( D => n1519, CK => CLK, Q => 
                           n14339, QN => n9482);
   REGISTERS_reg_26_16_inst : DFF_X1 port map( D => n1518, CK => CLK, Q => 
                           n14338, QN => n9483);
   REGISTERS_reg_26_15_inst : DFF_X1 port map( D => n1517, CK => CLK, Q => 
                           n14337, QN => n9484);
   REGISTERS_reg_26_14_inst : DFF_X1 port map( D => n1516, CK => CLK, Q => 
                           n14336, QN => n9485);
   REGISTERS_reg_26_13_inst : DFF_X1 port map( D => n1515, CK => CLK, Q => 
                           n14335, QN => n9486);
   REGISTERS_reg_26_12_inst : DFF_X1 port map( D => n1514, CK => CLK, Q => 
                           n14334, QN => n9487);
   REGISTERS_reg_26_11_inst : DFF_X1 port map( D => n1513, CK => CLK, Q => 
                           n14333, QN => n9488);
   REGISTERS_reg_26_10_inst : DFF_X1 port map( D => n1512, CK => CLK, Q => 
                           n14332, QN => n9489);
   REGISTERS_reg_26_9_inst : DFF_X1 port map( D => n1511, CK => CLK, Q => 
                           n14331, QN => n9490);
   REGISTERS_reg_26_8_inst : DFF_X1 port map( D => n1510, CK => CLK, Q => 
                           n14330, QN => n9491);
   REGISTERS_reg_26_7_inst : DFF_X1 port map( D => n1509, CK => CLK, Q => 
                           n14329, QN => n9492);
   REGISTERS_reg_26_6_inst : DFF_X1 port map( D => n1508, CK => CLK, Q => 
                           n14328, QN => n9493);
   REGISTERS_reg_26_5_inst : DFF_X1 port map( D => n1507, CK => CLK, Q => 
                           n14327, QN => n9494);
   REGISTERS_reg_26_4_inst : DFF_X1 port map( D => n1506, CK => CLK, Q => 
                           n14326, QN => n9495);
   REGISTERS_reg_26_3_inst : DFF_X1 port map( D => n1505, CK => CLK, Q => 
                           n14325, QN => n9496);
   REGISTERS_reg_26_2_inst : DFF_X1 port map( D => n1504, CK => CLK, Q => 
                           n14324, QN => n9497);
   REGISTERS_reg_26_1_inst : DFF_X1 port map( D => n1503, CK => CLK, Q => 
                           n14323, QN => n9498);
   REGISTERS_reg_26_0_inst : DFF_X1 port map( D => n1502, CK => CLK, Q => 
                           n14322, QN => n9499);
   REGISTERS_reg_27_31_inst : DFF_X1 port map( D => n1501, CK => CLK, Q => 
                           n_1448, QN => n9500);
   REGISTERS_reg_27_30_inst : DFF_X1 port map( D => n1500, CK => CLK, Q => 
                           n_1449, QN => n9501);
   REGISTERS_reg_27_29_inst : DFF_X1 port map( D => n1499, CK => CLK, Q => 
                           n_1450, QN => n9502);
   REGISTERS_reg_27_28_inst : DFF_X1 port map( D => n1498, CK => CLK, Q => 
                           n_1451, QN => n9503);
   REGISTERS_reg_27_27_inst : DFF_X1 port map( D => n1497, CK => CLK, Q => 
                           n_1452, QN => n9504);
   REGISTERS_reg_27_26_inst : DFF_X1 port map( D => n1496, CK => CLK, Q => 
                           n_1453, QN => n9505);
   REGISTERS_reg_27_25_inst : DFF_X1 port map( D => n1495, CK => CLK, Q => 
                           n_1454, QN => n9506);
   REGISTERS_reg_27_24_inst : DFF_X1 port map( D => n1494, CK => CLK, Q => 
                           n_1455, QN => n9507);
   REGISTERS_reg_27_23_inst : DFF_X1 port map( D => n1493, CK => CLK, Q => 
                           n_1456, QN => n9508);
   REGISTERS_reg_27_22_inst : DFF_X1 port map( D => n1492, CK => CLK, Q => 
                           n_1457, QN => n9509);
   REGISTERS_reg_27_21_inst : DFF_X1 port map( D => n1491, CK => CLK, Q => 
                           n_1458, QN => n9510);
   REGISTERS_reg_27_20_inst : DFF_X1 port map( D => n1490, CK => CLK, Q => 
                           n_1459, QN => n9511);
   REGISTERS_reg_27_19_inst : DFF_X1 port map( D => n1489, CK => CLK, Q => 
                           n_1460, QN => n9512);
   REGISTERS_reg_27_18_inst : DFF_X1 port map( D => n1488, CK => CLK, Q => 
                           n_1461, QN => n9513);
   REGISTERS_reg_27_17_inst : DFF_X1 port map( D => n1487, CK => CLK, Q => 
                           n_1462, QN => n9514);
   REGISTERS_reg_27_16_inst : DFF_X1 port map( D => n1486, CK => CLK, Q => 
                           n_1463, QN => n9515);
   REGISTERS_reg_27_15_inst : DFF_X1 port map( D => n1485, CK => CLK, Q => 
                           n_1464, QN => n9516);
   REGISTERS_reg_27_14_inst : DFF_X1 port map( D => n1484, CK => CLK, Q => 
                           n_1465, QN => n9517);
   REGISTERS_reg_27_13_inst : DFF_X1 port map( D => n1483, CK => CLK, Q => 
                           n_1466, QN => n9518);
   REGISTERS_reg_27_12_inst : DFF_X1 port map( D => n1482, CK => CLK, Q => 
                           n_1467, QN => n9519);
   REGISTERS_reg_27_11_inst : DFF_X1 port map( D => n1481, CK => CLK, Q => 
                           n_1468, QN => n9520);
   REGISTERS_reg_27_10_inst : DFF_X1 port map( D => n1480, CK => CLK, Q => 
                           n_1469, QN => n9521);
   REGISTERS_reg_27_9_inst : DFF_X1 port map( D => n1479, CK => CLK, Q => 
                           n_1470, QN => n9522);
   REGISTERS_reg_27_8_inst : DFF_X1 port map( D => n1478, CK => CLK, Q => 
                           n_1471, QN => n9523);
   REGISTERS_reg_27_7_inst : DFF_X1 port map( D => n1477, CK => CLK, Q => 
                           n_1472, QN => n9524);
   REGISTERS_reg_27_6_inst : DFF_X1 port map( D => n1476, CK => CLK, Q => 
                           n_1473, QN => n9525);
   REGISTERS_reg_27_5_inst : DFF_X1 port map( D => n1475, CK => CLK, Q => 
                           n_1474, QN => n9526);
   REGISTERS_reg_27_4_inst : DFF_X1 port map( D => n1474, CK => CLK, Q => 
                           n_1475, QN => n9527);
   REGISTERS_reg_27_3_inst : DFF_X1 port map( D => n1473, CK => CLK, Q => 
                           n_1476, QN => n9528);
   REGISTERS_reg_27_2_inst : DFF_X1 port map( D => n1472, CK => CLK, Q => 
                           n_1477, QN => n9529);
   REGISTERS_reg_27_1_inst : DFF_X1 port map( D => n1471, CK => CLK, Q => 
                           n_1478, QN => n9530);
   REGISTERS_reg_27_0_inst : DFF_X1 port map( D => n1470, CK => CLK, Q => 
                           n_1479, QN => n9531);
   REGISTERS_reg_28_31_inst : DFF_X1 port map( D => n1469, CK => CLK, Q => 
                           n14385, QN => n9532);
   REGISTERS_reg_28_30_inst : DFF_X1 port map( D => n1468, CK => CLK, Q => 
                           n14384, QN => n9533);
   REGISTERS_reg_28_29_inst : DFF_X1 port map( D => n1467, CK => CLK, Q => 
                           n14383, QN => n9534);
   REGISTERS_reg_28_28_inst : DFF_X1 port map( D => n1466, CK => CLK, Q => 
                           n14382, QN => n9535);
   REGISTERS_reg_28_27_inst : DFF_X1 port map( D => n1465, CK => CLK, Q => 
                           n14381, QN => n9536);
   REGISTERS_reg_28_26_inst : DFF_X1 port map( D => n1464, CK => CLK, Q => 
                           n14380, QN => n9537);
   REGISTERS_reg_28_25_inst : DFF_X1 port map( D => n1463, CK => CLK, Q => 
                           n14379, QN => n9538);
   REGISTERS_reg_28_24_inst : DFF_X1 port map( D => n1462, CK => CLK, Q => 
                           n14378, QN => n9539);
   REGISTERS_reg_28_23_inst : DFF_X1 port map( D => n1461, CK => CLK, Q => 
                           n14377, QN => n9540);
   REGISTERS_reg_28_22_inst : DFF_X1 port map( D => n1460, CK => CLK, Q => 
                           n14376, QN => n9541);
   REGISTERS_reg_28_21_inst : DFF_X1 port map( D => n1459, CK => CLK, Q => 
                           n14375, QN => n9542);
   REGISTERS_reg_28_20_inst : DFF_X1 port map( D => n1458, CK => CLK, Q => 
                           n14374, QN => n9543);
   REGISTERS_reg_28_19_inst : DFF_X1 port map( D => n1457, CK => CLK, Q => 
                           n14373, QN => n9544);
   REGISTERS_reg_28_18_inst : DFF_X1 port map( D => n1456, CK => CLK, Q => 
                           n14372, QN => n9545);
   REGISTERS_reg_28_17_inst : DFF_X1 port map( D => n1455, CK => CLK, Q => 
                           n14371, QN => n9546);
   REGISTERS_reg_28_16_inst : DFF_X1 port map( D => n1454, CK => CLK, Q => 
                           n14370, QN => n9547);
   REGISTERS_reg_28_15_inst : DFF_X1 port map( D => n1453, CK => CLK, Q => 
                           n14369, QN => n9548);
   REGISTERS_reg_28_14_inst : DFF_X1 port map( D => n1452, CK => CLK, Q => 
                           n14368, QN => n9549);
   REGISTERS_reg_28_13_inst : DFF_X1 port map( D => n1451, CK => CLK, Q => 
                           n14367, QN => n9550);
   REGISTERS_reg_28_12_inst : DFF_X1 port map( D => n1450, CK => CLK, Q => 
                           n14366, QN => n9551);
   REGISTERS_reg_28_11_inst : DFF_X1 port map( D => n1449, CK => CLK, Q => 
                           n14365, QN => n9552);
   REGISTERS_reg_28_10_inst : DFF_X1 port map( D => n1448, CK => CLK, Q => 
                           n14364, QN => n9553);
   REGISTERS_reg_28_9_inst : DFF_X1 port map( D => n1447, CK => CLK, Q => 
                           n14363, QN => n9554);
   REGISTERS_reg_28_8_inst : DFF_X1 port map( D => n1446, CK => CLK, Q => 
                           n14362, QN => n9555);
   REGISTERS_reg_28_7_inst : DFF_X1 port map( D => n1445, CK => CLK, Q => 
                           n14361, QN => n9556);
   REGISTERS_reg_28_6_inst : DFF_X1 port map( D => n1444, CK => CLK, Q => 
                           n14360, QN => n9557);
   REGISTERS_reg_28_5_inst : DFF_X1 port map( D => n1443, CK => CLK, Q => 
                           n14359, QN => n9558);
   REGISTERS_reg_28_4_inst : DFF_X1 port map( D => n1442, CK => CLK, Q => 
                           n14358, QN => n9559);
   REGISTERS_reg_28_3_inst : DFF_X1 port map( D => n1441, CK => CLK, Q => 
                           n14357, QN => n9560);
   REGISTERS_reg_28_2_inst : DFF_X1 port map( D => n1440, CK => CLK, Q => 
                           n14356, QN => n9561);
   REGISTERS_reg_28_1_inst : DFF_X1 port map( D => n1439, CK => CLK, Q => 
                           n14355, QN => n9562);
   REGISTERS_reg_28_0_inst : DFF_X1 port map( D => n1438, CK => CLK, Q => 
                           n14354, QN => n9563);
   REGISTERS_reg_29_31_inst : DFF_X1 port map( D => n1437, CK => CLK, Q => 
                           n13979, QN => n9564);
   REGISTERS_reg_29_30_inst : DFF_X1 port map( D => n1436, CK => CLK, Q => 
                           n13978, QN => n9565);
   REGISTERS_reg_29_29_inst : DFF_X1 port map( D => n1435, CK => CLK, Q => 
                           n13977, QN => n9566);
   REGISTERS_reg_29_28_inst : DFF_X1 port map( D => n1434, CK => CLK, Q => 
                           n13976, QN => n9567);
   REGISTERS_reg_29_27_inst : DFF_X1 port map( D => n1433, CK => CLK, Q => 
                           n13975, QN => n9568);
   REGISTERS_reg_29_26_inst : DFF_X1 port map( D => n1432, CK => CLK, Q => 
                           n13974, QN => n9569);
   REGISTERS_reg_29_25_inst : DFF_X1 port map( D => n1431, CK => CLK, Q => 
                           n13973, QN => n9570);
   REGISTERS_reg_29_24_inst : DFF_X1 port map( D => n1430, CK => CLK, Q => 
                           n13972, QN => n9571);
   REGISTERS_reg_29_23_inst : DFF_X1 port map( D => n1429, CK => CLK, Q => 
                           n13971, QN => n9572);
   REGISTERS_reg_29_22_inst : DFF_X1 port map( D => n1428, CK => CLK, Q => 
                           n13970, QN => n9573);
   REGISTERS_reg_29_21_inst : DFF_X1 port map( D => n1427, CK => CLK, Q => 
                           n13969, QN => n9574);
   REGISTERS_reg_29_20_inst : DFF_X1 port map( D => n1426, CK => CLK, Q => 
                           n13968, QN => n9575);
   REGISTERS_reg_29_19_inst : DFF_X1 port map( D => n1425, CK => CLK, Q => 
                           n13967, QN => n9576);
   REGISTERS_reg_29_18_inst : DFF_X1 port map( D => n1424, CK => CLK, Q => 
                           n13966, QN => n9577);
   REGISTERS_reg_29_17_inst : DFF_X1 port map( D => n1423, CK => CLK, Q => 
                           n13965, QN => n9578);
   REGISTERS_reg_29_16_inst : DFF_X1 port map( D => n1422, CK => CLK, Q => 
                           n13964, QN => n9579);
   REGISTERS_reg_29_15_inst : DFF_X1 port map( D => n1421, CK => CLK, Q => 
                           n13963, QN => n9580);
   REGISTERS_reg_29_14_inst : DFF_X1 port map( D => n1420, CK => CLK, Q => 
                           n13962, QN => n9581);
   REGISTERS_reg_29_13_inst : DFF_X1 port map( D => n1419, CK => CLK, Q => 
                           n13961, QN => n9582);
   REGISTERS_reg_29_12_inst : DFF_X1 port map( D => n1418, CK => CLK, Q => 
                           n13960, QN => n9583);
   REGISTERS_reg_29_11_inst : DFF_X1 port map( D => n1417, CK => CLK, Q => 
                           n13959, QN => n9584);
   REGISTERS_reg_29_10_inst : DFF_X1 port map( D => n1416, CK => CLK, Q => 
                           n13958, QN => n9585);
   REGISTERS_reg_29_9_inst : DFF_X1 port map( D => n1415, CK => CLK, Q => 
                           n13957, QN => n9586);
   REGISTERS_reg_29_8_inst : DFF_X1 port map( D => n1414, CK => CLK, Q => 
                           n13956, QN => n9587);
   REGISTERS_reg_29_7_inst : DFF_X1 port map( D => n1413, CK => CLK, Q => 
                           n13955, QN => n9588);
   REGISTERS_reg_29_6_inst : DFF_X1 port map( D => n1412, CK => CLK, Q => 
                           n13954, QN => n9589);
   REGISTERS_reg_29_5_inst : DFF_X1 port map( D => n1411, CK => CLK, Q => 
                           n13953, QN => n9590);
   REGISTERS_reg_29_4_inst : DFF_X1 port map( D => n1410, CK => CLK, Q => 
                           n13952, QN => n9591);
   REGISTERS_reg_29_3_inst : DFF_X1 port map( D => n1409, CK => CLK, Q => 
                           n13951, QN => n9592);
   REGISTERS_reg_29_2_inst : DFF_X1 port map( D => n1408, CK => CLK, Q => 
                           n13950, QN => n9593);
   REGISTERS_reg_29_1_inst : DFF_X1 port map( D => n1407, CK => CLK, Q => 
                           n13949, QN => n9594);
   REGISTERS_reg_29_0_inst : DFF_X1 port map( D => n1406, CK => CLK, Q => 
                           n13948, QN => n9595);
   REGISTERS_reg_30_31_inst : DFF_X1 port map( D => n1405, CK => CLK, Q => 
                           n_1480, QN => n9596);
   REGISTERS_reg_30_30_inst : DFF_X1 port map( D => n1404, CK => CLK, Q => 
                           n_1481, QN => n9597);
   REGISTERS_reg_30_29_inst : DFF_X1 port map( D => n1403, CK => CLK, Q => 
                           n_1482, QN => n9598);
   REGISTERS_reg_30_28_inst : DFF_X1 port map( D => n1402, CK => CLK, Q => 
                           n_1483, QN => n9599);
   REGISTERS_reg_30_27_inst : DFF_X1 port map( D => n1401, CK => CLK, Q => 
                           n_1484, QN => n9600);
   REGISTERS_reg_30_26_inst : DFF_X1 port map( D => n1400, CK => CLK, Q => 
                           n_1485, QN => n9601);
   REGISTERS_reg_30_25_inst : DFF_X1 port map( D => n1399, CK => CLK, Q => 
                           n_1486, QN => n9602);
   REGISTERS_reg_30_24_inst : DFF_X1 port map( D => n1398, CK => CLK, Q => 
                           n_1487, QN => n9603);
   REGISTERS_reg_30_23_inst : DFF_X1 port map( D => n1397, CK => CLK, Q => 
                           n_1488, QN => n9604);
   REGISTERS_reg_30_22_inst : DFF_X1 port map( D => n1396, CK => CLK, Q => 
                           n_1489, QN => n9605);
   REGISTERS_reg_30_21_inst : DFF_X1 port map( D => n1395, CK => CLK, Q => 
                           n_1490, QN => n9606);
   REGISTERS_reg_30_20_inst : DFF_X1 port map( D => n1394, CK => CLK, Q => 
                           n_1491, QN => n9607);
   REGISTERS_reg_30_19_inst : DFF_X1 port map( D => n1393, CK => CLK, Q => 
                           n_1492, QN => n9608);
   REGISTERS_reg_30_18_inst : DFF_X1 port map( D => n1392, CK => CLK, Q => 
                           n_1493, QN => n9609);
   REGISTERS_reg_30_17_inst : DFF_X1 port map( D => n1391, CK => CLK, Q => 
                           n_1494, QN => n9610);
   REGISTERS_reg_30_16_inst : DFF_X1 port map( D => n1390, CK => CLK, Q => 
                           n_1495, QN => n9611);
   REGISTERS_reg_30_15_inst : DFF_X1 port map( D => n1389, CK => CLK, Q => 
                           n_1496, QN => n9612);
   REGISTERS_reg_30_14_inst : DFF_X1 port map( D => n1388, CK => CLK, Q => 
                           n_1497, QN => n9613);
   REGISTERS_reg_30_13_inst : DFF_X1 port map( D => n1387, CK => CLK, Q => 
                           n_1498, QN => n9614);
   REGISTERS_reg_30_12_inst : DFF_X1 port map( D => n1386, CK => CLK, Q => 
                           n_1499, QN => n9615);
   REGISTERS_reg_30_11_inst : DFF_X1 port map( D => n1385, CK => CLK, Q => 
                           n_1500, QN => n9616);
   REGISTERS_reg_30_10_inst : DFF_X1 port map( D => n1384, CK => CLK, Q => 
                           n_1501, QN => n9617);
   REGISTERS_reg_30_9_inst : DFF_X1 port map( D => n1383, CK => CLK, Q => 
                           n_1502, QN => n9618);
   REGISTERS_reg_30_8_inst : DFF_X1 port map( D => n1382, CK => CLK, Q => 
                           n_1503, QN => n9619);
   REGISTERS_reg_30_7_inst : DFF_X1 port map( D => n1381, CK => CLK, Q => 
                           n_1504, QN => n9620);
   REGISTERS_reg_30_6_inst : DFF_X1 port map( D => n1380, CK => CLK, Q => 
                           n_1505, QN => n9621);
   REGISTERS_reg_30_5_inst : DFF_X1 port map( D => n1379, CK => CLK, Q => 
                           n_1506, QN => n9622);
   REGISTERS_reg_30_4_inst : DFF_X1 port map( D => n1378, CK => CLK, Q => 
                           n_1507, QN => n9623);
   REGISTERS_reg_30_3_inst : DFF_X1 port map( D => n1377, CK => CLK, Q => 
                           n_1508, QN => n9624);
   REGISTERS_reg_30_2_inst : DFF_X1 port map( D => n1376, CK => CLK, Q => 
                           n_1509, QN => n9625);
   REGISTERS_reg_30_1_inst : DFF_X1 port map( D => n1375, CK => CLK, Q => 
                           n_1510, QN => n9626);
   REGISTERS_reg_30_0_inst : DFF_X1 port map( D => n1374, CK => CLK, Q => 
                           n_1511, QN => n9627);
   REGISTERS_reg_31_31_inst : DFF_X1 port map( D => n1373, CK => CLK, Q => 
                           n_1512, QN => n13727);
   REGISTERS_reg_31_30_inst : DFF_X1 port map( D => n1372, CK => CLK, Q => 
                           n_1513, QN => n13636);
   REGISTERS_reg_31_29_inst : DFF_X1 port map( D => n1371, CK => CLK, Q => 
                           n_1514, QN => n9630);
   REGISTERS_reg_31_28_inst : DFF_X1 port map( D => n1370, CK => CLK, Q => 
                           n_1515, QN => n9631);
   REGISTERS_reg_31_27_inst : DFF_X1 port map( D => n1369, CK => CLK, Q => 
                           n_1516, QN => n9632);
   REGISTERS_reg_31_26_inst : DFF_X1 port map( D => n1368, CK => CLK, Q => 
                           n_1517, QN => n9633);
   REGISTERS_reg_31_25_inst : DFF_X1 port map( D => n1367, CK => CLK, Q => 
                           n_1518, QN => n9634);
   REGISTERS_reg_31_24_inst : DFF_X1 port map( D => n1366, CK => CLK, Q => 
                           n_1519, QN => n9635);
   REGISTERS_reg_31_23_inst : DFF_X1 port map( D => n1365, CK => CLK, Q => 
                           n_1520, QN => n9636);
   REGISTERS_reg_31_22_inst : DFF_X1 port map( D => n1364, CK => CLK, Q => 
                           n_1521, QN => n9637);
   REGISTERS_reg_31_21_inst : DFF_X1 port map( D => n1363, CK => CLK, Q => 
                           n_1522, QN => n9638);
   REGISTERS_reg_31_20_inst : DFF_X1 port map( D => n1362, CK => CLK, Q => 
                           n_1523, QN => n9639);
   REGISTERS_reg_31_19_inst : DFF_X1 port map( D => n1361, CK => CLK, Q => 
                           n_1524, QN => n9640);
   REGISTERS_reg_31_18_inst : DFF_X1 port map( D => n1360, CK => CLK, Q => 
                           n_1525, QN => n9641);
   REGISTERS_reg_31_17_inst : DFF_X1 port map( D => n1359, CK => CLK, Q => 
                           n_1526, QN => n9642);
   REGISTERS_reg_31_16_inst : DFF_X1 port map( D => n1358, CK => CLK, Q => 
                           n_1527, QN => n9643);
   REGISTERS_reg_31_15_inst : DFF_X1 port map( D => n1357, CK => CLK, Q => 
                           n_1528, QN => n9644);
   REGISTERS_reg_31_14_inst : DFF_X1 port map( D => n1356, CK => CLK, Q => 
                           n_1529, QN => n9645);
   REGISTERS_reg_31_13_inst : DFF_X1 port map( D => n1355, CK => CLK, Q => 
                           n_1530, QN => n9646);
   REGISTERS_reg_31_12_inst : DFF_X1 port map( D => n1354, CK => CLK, Q => 
                           n_1531, QN => n9647);
   REGISTERS_reg_31_11_inst : DFF_X1 port map( D => n1353, CK => CLK, Q => 
                           n_1532, QN => n9648);
   REGISTERS_reg_31_10_inst : DFF_X1 port map( D => n1352, CK => CLK, Q => 
                           n_1533, QN => n13726);
   REGISTERS_reg_31_9_inst : DFF_X1 port map( D => n1351, CK => CLK, Q => 
                           n_1534, QN => n13725);
   REGISTERS_reg_31_8_inst : DFF_X1 port map( D => n1350, CK => CLK, Q => 
                           n_1535, QN => n13724);
   REGISTERS_reg_31_7_inst : DFF_X1 port map( D => n1349, CK => CLK, Q => 
                           n_1536, QN => n13643);
   REGISTERS_reg_31_6_inst : DFF_X1 port map( D => n1348, CK => CLK, Q => 
                           n_1537, QN => n13642);
   REGISTERS_reg_31_5_inst : DFF_X1 port map( D => n1347, CK => CLK, Q => 
                           n_1538, QN => n13641);
   REGISTERS_reg_31_4_inst : DFF_X1 port map( D => n1346, CK => CLK, Q => 
                           n_1539, QN => n13640);
   REGISTERS_reg_31_3_inst : DFF_X1 port map( D => n1345, CK => CLK, Q => 
                           n_1540, QN => n13639);
   REGISTERS_reg_31_2_inst : DFF_X1 port map( D => n1344, CK => CLK, Q => 
                           n_1541, QN => n13638);
   REGISTERS_reg_31_1_inst : DFF_X1 port map( D => n1343, CK => CLK, Q => 
                           n_1542, QN => n13637);
   REGISTERS_reg_31_0_inst : DFF_X1 port map( D => n1342, CK => CLK, Q => 
                           n_1543, QN => n9659);
   OUT1_reg_31_inst : DFF_X1 port map( D => n1341, CK => CLK, Q => OUT1(31), QN
                           => n13191);
   OUT1_reg_30_inst : DFF_X1 port map( D => n1340, CK => CLK, Q => OUT1(30), QN
                           => n13190);
   OUT1_reg_29_inst : DFF_X1 port map( D => n1339, CK => CLK, Q => OUT1(29), QN
                           => n13251);
   OUT1_reg_28_inst : DFF_X1 port map( D => n1338, CK => CLK, Q => OUT1(28), QN
                           => n13250);
   OUT1_reg_27_inst : DFF_X1 port map( D => n1337, CK => CLK, Q => OUT1(27), QN
                           => n13249);
   OUT1_reg_26_inst : DFF_X1 port map( D => n1336, CK => CLK, Q => OUT1(26), QN
                           => n13248);
   OUT1_reg_25_inst : DFF_X1 port map( D => n1335, CK => CLK, Q => OUT1(25), QN
                           => n13247);
   OUT1_reg_24_inst : DFF_X1 port map( D => n1334, CK => CLK, Q => OUT1(24), QN
                           => n13246);
   OUT1_reg_23_inst : DFF_X1 port map( D => n1333, CK => CLK, Q => OUT1(23), QN
                           => n13245);
   OUT1_reg_22_inst : DFF_X1 port map( D => n1332, CK => CLK, Q => OUT1(22), QN
                           => n13244);
   OUT1_reg_21_inst : DFF_X1 port map( D => n1331, CK => CLK, Q => OUT1(21), QN
                           => n13243);
   OUT1_reg_20_inst : DFF_X1 port map( D => n1330, CK => CLK, Q => OUT1(20), QN
                           => n13242);
   OUT1_reg_19_inst : DFF_X1 port map( D => n1329, CK => CLK, Q => OUT1(19), QN
                           => n13241);
   OUT1_reg_18_inst : DFF_X1 port map( D => n1328, CK => CLK, Q => OUT1(18), QN
                           => n13240);
   OUT1_reg_17_inst : DFF_X1 port map( D => n1327, CK => CLK, Q => OUT1(17), QN
                           => n13239);
   OUT1_reg_16_inst : DFF_X1 port map( D => n1326, CK => CLK, Q => OUT1(16), QN
                           => n13238);
   OUT1_reg_15_inst : DFF_X1 port map( D => n1325, CK => CLK, Q => OUT1(15), QN
                           => n13237);
   OUT1_reg_14_inst : DFF_X1 port map( D => n1324, CK => CLK, Q => OUT1(14), QN
                           => n13236);
   OUT1_reg_13_inst : DFF_X1 port map( D => n1323, CK => CLK, Q => OUT1(13), QN
                           => n13235);
   OUT1_reg_12_inst : DFF_X1 port map( D => n1322, CK => CLK, Q => OUT1(12), QN
                           => n13234);
   OUT1_reg_11_inst : DFF_X1 port map( D => n1321, CK => CLK, Q => OUT1(11), QN
                           => n13233);
   OUT1_reg_10_inst : DFF_X1 port map( D => n1320, CK => CLK, Q => OUT1(10), QN
                           => n13232);
   OUT1_reg_9_inst : DFF_X1 port map( D => n1319, CK => CLK, Q => OUT1(9), QN 
                           => n13231);
   OUT1_reg_8_inst : DFF_X1 port map( D => n1318, CK => CLK, Q => OUT1(8), QN 
                           => n13230);
   OUT1_reg_7_inst : DFF_X1 port map( D => n1317, CK => CLK, Q => OUT1(7), QN 
                           => n13229);
   OUT1_reg_6_inst : DFF_X1 port map( D => n1316, CK => CLK, Q => OUT1(6), QN 
                           => n13228);
   OUT1_reg_5_inst : DFF_X1 port map( D => n1315, CK => CLK, Q => OUT1(5), QN 
                           => n13227);
   OUT1_reg_4_inst : DFF_X1 port map( D => n1314, CK => CLK, Q => OUT1(4), QN 
                           => n13226);
   OUT1_reg_3_inst : DFF_X1 port map( D => n1313, CK => CLK, Q => OUT1(3), QN 
                           => n13225);
   OUT1_reg_2_inst : DFF_X1 port map( D => n1312, CK => CLK, Q => OUT1(2), QN 
                           => n13224);
   OUT1_reg_1_inst : DFF_X1 port map( D => n1311, CK => CLK, Q => OUT1(1), QN 
                           => n13223);
   OUT1_reg_0_inst : DFF_X1 port map( D => n1310, CK => CLK, Q => OUT1(0), QN 
                           => n13222);
   OUT2_reg_31_inst : DFF_X1 port map( D => n1309, CK => CLK, Q => OUT2(31), QN
                           => n13189);
   OUT2_reg_30_inst : DFF_X1 port map( D => n1308, CK => CLK, Q => OUT2(30), QN
                           => n13188);
   OUT2_reg_29_inst : DFF_X1 port map( D => n1307, CK => CLK, Q => OUT2(29), QN
                           => n13221);
   OUT2_reg_28_inst : DFF_X1 port map( D => n1306, CK => CLK, Q => OUT2(28), QN
                           => n13220);
   OUT2_reg_27_inst : DFF_X1 port map( D => n1305, CK => CLK, Q => OUT2(27), QN
                           => n13219);
   OUT2_reg_26_inst : DFF_X1 port map( D => n1304, CK => CLK, Q => OUT2(26), QN
                           => n13218);
   OUT2_reg_25_inst : DFF_X1 port map( D => n1303, CK => CLK, Q => OUT2(25), QN
                           => n13217);
   OUT2_reg_24_inst : DFF_X1 port map( D => n1302, CK => CLK, Q => OUT2(24), QN
                           => n13216);
   OUT2_reg_23_inst : DFF_X1 port map( D => n1301, CK => CLK, Q => OUT2(23), QN
                           => n13215);
   OUT2_reg_22_inst : DFF_X1 port map( D => n1300, CK => CLK, Q => OUT2(22), QN
                           => n13214);
   OUT2_reg_21_inst : DFF_X1 port map( D => n1299, CK => CLK, Q => OUT2(21), QN
                           => n13213);
   OUT2_reg_20_inst : DFF_X1 port map( D => n1298, CK => CLK, Q => OUT2(20), QN
                           => n13212);
   OUT2_reg_19_inst : DFF_X1 port map( D => n1297, CK => CLK, Q => OUT2(19), QN
                           => n13211);
   OUT2_reg_18_inst : DFF_X1 port map( D => n1296, CK => CLK, Q => OUT2(18), QN
                           => n13210);
   OUT2_reg_17_inst : DFF_X1 port map( D => n1295, CK => CLK, Q => OUT2(17), QN
                           => n13209);
   OUT2_reg_16_inst : DFF_X1 port map( D => n1294, CK => CLK, Q => OUT2(16), QN
                           => n13208);
   OUT2_reg_15_inst : DFF_X1 port map( D => n1293, CK => CLK, Q => OUT2(15), QN
                           => n13207);
   OUT2_reg_14_inst : DFF_X1 port map( D => n1292, CK => CLK, Q => OUT2(14), QN
                           => n13206);
   OUT2_reg_13_inst : DFF_X1 port map( D => n1291, CK => CLK, Q => OUT2(13), QN
                           => n13205);
   OUT2_reg_12_inst : DFF_X1 port map( D => n1290, CK => CLK, Q => OUT2(12), QN
                           => n13204);
   OUT2_reg_11_inst : DFF_X1 port map( D => n1289, CK => CLK, Q => OUT2(11), QN
                           => n13203);
   OUT2_reg_10_inst : DFF_X1 port map( D => n1288, CK => CLK, Q => OUT2(10), QN
                           => n13202);
   OUT2_reg_9_inst : DFF_X1 port map( D => n1287, CK => CLK, Q => OUT2(9), QN 
                           => n13201);
   OUT2_reg_8_inst : DFF_X1 port map( D => n1286, CK => CLK, Q => OUT2(8), QN 
                           => n13200);
   OUT2_reg_7_inst : DFF_X1 port map( D => n1285, CK => CLK, Q => OUT2(7), QN 
                           => n13199);
   OUT2_reg_6_inst : DFF_X1 port map( D => n1284, CK => CLK, Q => OUT2(6), QN 
                           => n13198);
   OUT2_reg_5_inst : DFF_X1 port map( D => n1283, CK => CLK, Q => OUT2(5), QN 
                           => n13197);
   OUT2_reg_4_inst : DFF_X1 port map( D => n1282, CK => CLK, Q => OUT2(4), QN 
                           => n13196);
   OUT2_reg_3_inst : DFF_X1 port map( D => n1281, CK => CLK, Q => OUT2(3), QN 
                           => n13195);
   OUT2_reg_2_inst : DFF_X1 port map( D => n1280, CK => CLK, Q => OUT2(2), QN 
                           => n13194);
   OUT2_reg_1_inst : DFF_X1 port map( D => n1279, CK => CLK, Q => OUT2(1), QN 
                           => n13193);
   OUT2_reg_0_inst : DFF_X1 port map( D => n1278, CK => CLK, Q => OUT2(0), QN 
                           => n13192);
   U9878 : NAND3_X1 port map( A1 => n10989, A2 => n10988, A3 => n11989, ZN => 
                           n11981);
   U9879 : NAND3_X1 port map( A1 => n11989, A2 => n10988, A3 => ADD_WR(2), ZN 
                           => n11991);
   U9880 : NAND3_X1 port map( A1 => n11989, A2 => n10989, A3 => ADD_WR(3), ZN 
                           => n11996);
   U9881 : NAND3_X1 port map( A1 => ADD_WR(2), A2 => n11989, A3 => ADD_WR(3), 
                           ZN => n12001);
   U9882 : NAND3_X1 port map( A1 => n10989, A2 => n10988, A3 => n12010, ZN => 
                           n12006);
   U9883 : NAND3_X1 port map( A1 => ADD_WR(2), A2 => n10988, A3 => n12010, ZN 
                           => n12012);
   U9884 : NAND3_X1 port map( A1 => ADD_WR(3), A2 => n10989, A3 => n12010, ZN 
                           => n12017);
   U9885 : NAND3_X1 port map( A1 => ADD_WR(3), A2 => ADD_WR(2), A3 => n12010, 
                           ZN => n12022);
   U9894 : AND3_X1 port map( A1 => ADD_RD2(3), A2 => n11005, A3 => ADD_RD2(4), 
                           ZN => n14044);
   U9895 : AND3_X1 port map( A1 => ADD_RD1(3), A2 => n10997, A3 => ADD_RD1(4), 
                           ZN => n14045);
   U9896 : INV_X1 port map( A => n14924, ZN => n14917);
   U9897 : INV_X1 port map( A => n15161, ZN => n15154);
   U9898 : INV_X1 port map( A => n14798, ZN => n14791);
   U9899 : INV_X1 port map( A => n14807, ZN => n14800);
   U9900 : INV_X1 port map( A => n14816, ZN => n14809);
   U9901 : INV_X1 port map( A => n14825, ZN => n14818);
   U9902 : INV_X1 port map( A => n14834, ZN => n14827);
   U9903 : INV_X1 port map( A => n14843, ZN => n14836);
   U9904 : INV_X1 port map( A => n14852, ZN => n14845);
   U9905 : INV_X1 port map( A => n14933, ZN => n14926);
   U9906 : INV_X1 port map( A => n14969, ZN => n14962);
   U9907 : INV_X1 port map( A => n14861, ZN => n14854);
   U9908 : INV_X1 port map( A => n14870, ZN => n14863);
   U9909 : INV_X1 port map( A => n14879, ZN => n14872);
   U9910 : INV_X1 port map( A => n14888, ZN => n14881);
   U9911 : INV_X1 port map( A => n14897, ZN => n14890);
   U9912 : INV_X1 port map( A => n14906, ZN => n14899);
   U9913 : INV_X1 port map( A => n14915, ZN => n14908);
   U9914 : INV_X1 port map( A => n14942, ZN => n14935);
   U9915 : INV_X1 port map( A => n14951, ZN => n14944);
   U9916 : INV_X1 port map( A => n14960, ZN => n14953);
   U9917 : INV_X1 port map( A => n14978, ZN => n14971);
   U9918 : INV_X1 port map( A => n14987, ZN => n14980);
   U9919 : INV_X1 port map( A => n14996, ZN => n14989);
   U9920 : INV_X1 port map( A => n15005, ZN => n14998);
   U9921 : INV_X1 port map( A => n15014, ZN => n15007);
   U9922 : INV_X1 port map( A => n15023, ZN => n15016);
   U9923 : INV_X1 port map( A => n15032, ZN => n15025);
   U9924 : INV_X1 port map( A => n15041, ZN => n15034);
   U9925 : INV_X1 port map( A => n15050, ZN => n15043);
   U9926 : INV_X1 port map( A => n15059, ZN => n15052);
   U9927 : BUF_X1 port map( A => n12640, Z => n14626);
   U9928 : BUF_X1 port map( A => n12640, Z => n14627);
   U9929 : BUF_X1 port map( A => n12059, Z => n14724);
   U9930 : BUF_X1 port map( A => n12059, Z => n14725);
   U9931 : BUF_X1 port map( A => n12633, Z => n14644);
   U9932 : BUF_X1 port map( A => n12633, Z => n14645);
   U9933 : BUF_X1 port map( A => n12052, Z => n14742);
   U9934 : BUF_X1 port map( A => n12052, Z => n14743);
   U9935 : BUF_X1 port map( A => n12636, Z => n14635);
   U9936 : BUF_X1 port map( A => n12636, Z => n14636);
   U9937 : BUF_X1 port map( A => n12055, Z => n14733);
   U9938 : BUF_X1 port map( A => n12055, Z => n14734);
   U9939 : BUF_X1 port map( A => n12653, Z => n14597);
   U9940 : BUF_X1 port map( A => n12656, Z => n14588);
   U9941 : BUF_X1 port map( A => n12653, Z => n14596);
   U9942 : BUF_X1 port map( A => n12656, Z => n14587);
   U9943 : BUF_X1 port map( A => n12072, Z => n14695);
   U9944 : BUF_X1 port map( A => n12075, Z => n14686);
   U9945 : BUF_X1 port map( A => n12072, Z => n14694);
   U9946 : BUF_X1 port map( A => n12075, Z => n14685);
   U9947 : BUF_X1 port map( A => n12640, Z => n14628);
   U9948 : BUF_X1 port map( A => n12059, Z => n14726);
   U9949 : BUF_X1 port map( A => n12633, Z => n14646);
   U9950 : BUF_X1 port map( A => n12052, Z => n14744);
   U9951 : BUF_X1 port map( A => n12636, Z => n14637);
   U9952 : BUF_X1 port map( A => n12055, Z => n14735);
   U9953 : BUF_X1 port map( A => n12653, Z => n14598);
   U9954 : BUF_X1 port map( A => n12656, Z => n14589);
   U9955 : BUF_X1 port map( A => n12072, Z => n14696);
   U9956 : BUF_X1 port map( A => n12075, Z => n14687);
   U9957 : BUF_X1 port map( A => n14925, Z => n14918);
   U9958 : BUF_X1 port map( A => n14925, Z => n14919);
   U9959 : BUF_X1 port map( A => n14925, Z => n14920);
   U9960 : BUF_X1 port map( A => n14925, Z => n14921);
   U9961 : BUF_X1 port map( A => n14925, Z => n14922);
   U9962 : BUF_X1 port map( A => n14925, Z => n14923);
   U9963 : BUF_X1 port map( A => n15162, Z => n15155);
   U9964 : BUF_X1 port map( A => n15162, Z => n15156);
   U9965 : BUF_X1 port map( A => n15162, Z => n15157);
   U9966 : BUF_X1 port map( A => n15162, Z => n15158);
   U9967 : BUF_X1 port map( A => n15162, Z => n15159);
   U9968 : BUF_X1 port map( A => n15162, Z => n15160);
   U9969 : BUF_X1 port map( A => n14925, Z => n14924);
   U9970 : BUF_X1 port map( A => n15162, Z => n15161);
   U9971 : BUF_X1 port map( A => n14790, Z => n14781);
   U9972 : BUF_X1 port map( A => n14790, Z => n14782);
   U9973 : BUF_X1 port map( A => n14790, Z => n14783);
   U9974 : BUF_X1 port map( A => n14790, Z => n14784);
   U9975 : BUF_X1 port map( A => n14789, Z => n14785);
   U9976 : BUF_X1 port map( A => n14787, Z => n14786);
   U9977 : BUF_X1 port map( A => n14790, Z => n14787);
   U9978 : BUF_X1 port map( A => n14789, Z => n14788);
   U9979 : BUF_X1 port map( A => n14790, Z => n14789);
   U9980 : INV_X1 port map( A => n14044, ZN => n14671);
   U9981 : INV_X1 port map( A => n14044, ZN => n14672);
   U9982 : INV_X1 port map( A => n14045, ZN => n14769);
   U9983 : INV_X1 port map( A => n14045, ZN => n14770);
   U9984 : BUF_X1 port map( A => n12645, Z => n14617);
   U9985 : BUF_X1 port map( A => n12645, Z => n14618);
   U9986 : BUF_X1 port map( A => n12064, Z => n14715);
   U9987 : BUF_X1 port map( A => n12064, Z => n14716);
   U9988 : BUF_X1 port map( A => n12646, Z => n14614);
   U9989 : BUF_X1 port map( A => n12646, Z => n14615);
   U9990 : BUF_X1 port map( A => n12065, Z => n14712);
   U9991 : BUF_X1 port map( A => n12065, Z => n14713);
   U9992 : BUF_X1 port map( A => n12638, Z => n14629);
   U9993 : BUF_X1 port map( A => n12648, Z => n14608);
   U9994 : BUF_X1 port map( A => n12638, Z => n14630);
   U9995 : BUF_X1 port map( A => n12648, Z => n14609);
   U9996 : BUF_X1 port map( A => n12057, Z => n14727);
   U9997 : BUF_X1 port map( A => n12067, Z => n14706);
   U9998 : BUF_X1 port map( A => n12057, Z => n14728);
   U9999 : BUF_X1 port map( A => n12067, Z => n14707);
   U10000 : BUF_X1 port map( A => n12642, Z => n14620);
   U10001 : BUF_X1 port map( A => n12642, Z => n14621);
   U10002 : BUF_X1 port map( A => n12061, Z => n14718);
   U10003 : BUF_X1 port map( A => n12061, Z => n14719);
   U10004 : BUF_X1 port map( A => n12652, Z => n14599);
   U10005 : BUF_X1 port map( A => n12655, Z => n14590);
   U10006 : BUF_X1 port map( A => n12652, Z => n14600);
   U10007 : BUF_X1 port map( A => n12655, Z => n14591);
   U10008 : BUF_X1 port map( A => n12071, Z => n14697);
   U10009 : BUF_X1 port map( A => n12074, Z => n14688);
   U10010 : BUF_X1 port map( A => n12071, Z => n14698);
   U10011 : BUF_X1 port map( A => n12074, Z => n14689);
   U10012 : BUF_X1 port map( A => n12650, Z => n14605);
   U10013 : BUF_X1 port map( A => n12650, Z => n14606);
   U10014 : BUF_X1 port map( A => n12069, Z => n14703);
   U10015 : BUF_X1 port map( A => n12069, Z => n14704);
   U10016 : BUF_X1 port map( A => n12615, Z => n14679);
   U10017 : BUF_X1 port map( A => n12615, Z => n14680);
   U10018 : BUF_X1 port map( A => n12034, Z => n14777);
   U10019 : BUF_X1 port map( A => n12034, Z => n14778);
   U10020 : BUF_X1 port map( A => n12637, Z => n14632);
   U10021 : BUF_X1 port map( A => n12647, Z => n14611);
   U10022 : BUF_X1 port map( A => n12637, Z => n14633);
   U10023 : BUF_X1 port map( A => n12647, Z => n14612);
   U10024 : BUF_X1 port map( A => n12056, Z => n14730);
   U10025 : BUF_X1 port map( A => n12066, Z => n14709);
   U10026 : BUF_X1 port map( A => n12056, Z => n14731);
   U10027 : BUF_X1 port map( A => n12066, Z => n14710);
   U10028 : BUF_X1 port map( A => n12645, Z => n14619);
   U10029 : BUF_X1 port map( A => n12064, Z => n14717);
   U10030 : BUF_X1 port map( A => n12631, Z => n14650);
   U10031 : BUF_X1 port map( A => n12631, Z => n14651);
   U10032 : BUF_X1 port map( A => n12050, Z => n14748);
   U10033 : BUF_X1 port map( A => n12050, Z => n14749);
   U10034 : BUF_X1 port map( A => n12634, Z => n14641);
   U10035 : BUF_X1 port map( A => n12634, Z => n14642);
   U10036 : BUF_X1 port map( A => n12053, Z => n14739);
   U10037 : BUF_X1 port map( A => n12053, Z => n14740);
   U10038 : BUF_X1 port map( A => n12632, Z => n14647);
   U10039 : BUF_X1 port map( A => n12632, Z => n14648);
   U10040 : BUF_X1 port map( A => n12051, Z => n14745);
   U10041 : BUF_X1 port map( A => n12051, Z => n14746);
   U10042 : BUF_X1 port map( A => n12635, Z => n14638);
   U10043 : BUF_X1 port map( A => n12635, Z => n14639);
   U10044 : BUF_X1 port map( A => n12054, Z => n14736);
   U10045 : BUF_X1 port map( A => n12054, Z => n14737);
   U10046 : BUF_X1 port map( A => n12646, Z => n14616);
   U10047 : BUF_X1 port map( A => n12065, Z => n14714);
   U10048 : BUF_X1 port map( A => n12641, Z => n14624);
   U10049 : BUF_X1 port map( A => n12651, Z => n14603);
   U10050 : BUF_X1 port map( A => n12641, Z => n14623);
   U10051 : BUF_X1 port map( A => n12651, Z => n14602);
   U10052 : BUF_X1 port map( A => n12060, Z => n14722);
   U10053 : BUF_X1 port map( A => n12070, Z => n14701);
   U10054 : BUF_X1 port map( A => n12060, Z => n14721);
   U10055 : BUF_X1 port map( A => n12070, Z => n14700);
   U10056 : BUF_X1 port map( A => n12654, Z => n14594);
   U10057 : BUF_X1 port map( A => n12657, Z => n14585);
   U10058 : BUF_X1 port map( A => n12654, Z => n14593);
   U10059 : BUF_X1 port map( A => n12657, Z => n14584);
   U10060 : BUF_X1 port map( A => n12073, Z => n14692);
   U10061 : BUF_X1 port map( A => n12076, Z => n14683);
   U10062 : BUF_X1 port map( A => n12073, Z => n14691);
   U10063 : BUF_X1 port map( A => n12076, Z => n14682);
   U10064 : BUF_X1 port map( A => n12638, Z => n14631);
   U10065 : BUF_X1 port map( A => n12648, Z => n14610);
   U10066 : BUF_X1 port map( A => n12057, Z => n14729);
   U10067 : BUF_X1 port map( A => n12067, Z => n14708);
   U10068 : BUF_X1 port map( A => n12642, Z => n14622);
   U10069 : BUF_X1 port map( A => n12061, Z => n14720);
   U10070 : BUF_X1 port map( A => n12652, Z => n14601);
   U10071 : BUF_X1 port map( A => n12655, Z => n14592);
   U10072 : BUF_X1 port map( A => n12071, Z => n14699);
   U10073 : BUF_X1 port map( A => n12074, Z => n14690);
   U10074 : BUF_X1 port map( A => n12650, Z => n14607);
   U10075 : BUF_X1 port map( A => n12069, Z => n14705);
   U10076 : BUF_X1 port map( A => n12615, Z => n14681);
   U10077 : BUF_X1 port map( A => n12034, Z => n14779);
   U10078 : BUF_X1 port map( A => n12637, Z => n14634);
   U10079 : BUF_X1 port map( A => n12647, Z => n14613);
   U10080 : BUF_X1 port map( A => n12056, Z => n14732);
   U10081 : BUF_X1 port map( A => n12066, Z => n14711);
   U10082 : BUF_X1 port map( A => n12631, Z => n14652);
   U10083 : BUF_X1 port map( A => n12050, Z => n14750);
   U10084 : BUF_X1 port map( A => n12634, Z => n14643);
   U10085 : BUF_X1 port map( A => n12053, Z => n14741);
   U10086 : BUF_X1 port map( A => n12632, Z => n14649);
   U10087 : BUF_X1 port map( A => n12051, Z => n14747);
   U10088 : BUF_X1 port map( A => n12635, Z => n14640);
   U10089 : BUF_X1 port map( A => n12054, Z => n14738);
   U10090 : BUF_X1 port map( A => n12641, Z => n14625);
   U10091 : BUF_X1 port map( A => n12651, Z => n14604);
   U10092 : BUF_X1 port map( A => n12060, Z => n14723);
   U10093 : BUF_X1 port map( A => n12070, Z => n14702);
   U10094 : BUF_X1 port map( A => n12654, Z => n14595);
   U10095 : BUF_X1 port map( A => n12657, Z => n14586);
   U10096 : BUF_X1 port map( A => n12073, Z => n14693);
   U10097 : BUF_X1 port map( A => n12076, Z => n14684);
   U10098 : NAND2_X1 port map( A1 => n14663, A2 => n13182, ZN => n12633);
   U10099 : NAND2_X1 port map( A1 => n14761, A2 => n12601, ZN => n12052);
   U10100 : NAND2_X1 port map( A1 => n14668, A2 => n13182, ZN => n12636);
   U10101 : NAND2_X1 port map( A1 => n14766, A2 => n12601, ZN => n12055);
   U10102 : BUF_X1 port map( A => n14799, Z => n14792);
   U10103 : BUF_X1 port map( A => n14799, Z => n14793);
   U10104 : BUF_X1 port map( A => n14799, Z => n14794);
   U10105 : BUF_X1 port map( A => n14799, Z => n14795);
   U10106 : BUF_X1 port map( A => n14799, Z => n14796);
   U10107 : BUF_X1 port map( A => n14799, Z => n14797);
   U10108 : BUF_X1 port map( A => n14808, Z => n14801);
   U10109 : BUF_X1 port map( A => n14808, Z => n14802);
   U10110 : BUF_X1 port map( A => n14808, Z => n14803);
   U10111 : BUF_X1 port map( A => n14808, Z => n14804);
   U10112 : BUF_X1 port map( A => n14808, Z => n14805);
   U10113 : BUF_X1 port map( A => n14808, Z => n14806);
   U10114 : BUF_X1 port map( A => n14817, Z => n14810);
   U10115 : BUF_X1 port map( A => n14817, Z => n14811);
   U10116 : BUF_X1 port map( A => n14817, Z => n14812);
   U10117 : BUF_X1 port map( A => n14817, Z => n14813);
   U10118 : BUF_X1 port map( A => n14817, Z => n14814);
   U10119 : BUF_X1 port map( A => n14817, Z => n14815);
   U10120 : BUF_X1 port map( A => n14826, Z => n14819);
   U10121 : BUF_X1 port map( A => n14826, Z => n14820);
   U10122 : BUF_X1 port map( A => n14826, Z => n14821);
   U10123 : BUF_X1 port map( A => n14826, Z => n14822);
   U10124 : BUF_X1 port map( A => n14826, Z => n14823);
   U10125 : BUF_X1 port map( A => n14826, Z => n14824);
   U10126 : BUF_X1 port map( A => n14835, Z => n14828);
   U10127 : BUF_X1 port map( A => n14835, Z => n14829);
   U10128 : BUF_X1 port map( A => n14835, Z => n14830);
   U10129 : BUF_X1 port map( A => n14835, Z => n14831);
   U10130 : BUF_X1 port map( A => n14835, Z => n14832);
   U10131 : BUF_X1 port map( A => n14835, Z => n14833);
   U10132 : BUF_X1 port map( A => n14844, Z => n14837);
   U10133 : BUF_X1 port map( A => n14844, Z => n14838);
   U10134 : BUF_X1 port map( A => n14844, Z => n14839);
   U10135 : BUF_X1 port map( A => n14844, Z => n14840);
   U10136 : BUF_X1 port map( A => n14844, Z => n14841);
   U10137 : BUF_X1 port map( A => n14844, Z => n14842);
   U10138 : BUF_X1 port map( A => n14853, Z => n14846);
   U10139 : BUF_X1 port map( A => n14853, Z => n14847);
   U10140 : BUF_X1 port map( A => n14853, Z => n14848);
   U10141 : BUF_X1 port map( A => n14853, Z => n14849);
   U10142 : BUF_X1 port map( A => n14853, Z => n14850);
   U10143 : BUF_X1 port map( A => n14853, Z => n14851);
   U10144 : BUF_X1 port map( A => n14862, Z => n14855);
   U10145 : BUF_X1 port map( A => n14862, Z => n14856);
   U10146 : BUF_X1 port map( A => n14862, Z => n14857);
   U10147 : BUF_X1 port map( A => n14862, Z => n14858);
   U10148 : BUF_X1 port map( A => n14862, Z => n14859);
   U10149 : BUF_X1 port map( A => n14862, Z => n14860);
   U10150 : BUF_X1 port map( A => n14871, Z => n14864);
   U10151 : BUF_X1 port map( A => n14871, Z => n14865);
   U10152 : BUF_X1 port map( A => n14871, Z => n14866);
   U10153 : BUF_X1 port map( A => n14871, Z => n14867);
   U10154 : BUF_X1 port map( A => n14871, Z => n14868);
   U10155 : BUF_X1 port map( A => n14871, Z => n14869);
   U10156 : BUF_X1 port map( A => n14880, Z => n14873);
   U10157 : BUF_X1 port map( A => n14880, Z => n14874);
   U10158 : BUF_X1 port map( A => n14880, Z => n14875);
   U10159 : BUF_X1 port map( A => n14880, Z => n14876);
   U10160 : BUF_X1 port map( A => n14880, Z => n14877);
   U10161 : BUF_X1 port map( A => n14880, Z => n14878);
   U10162 : BUF_X1 port map( A => n14889, Z => n14882);
   U10163 : BUF_X1 port map( A => n14889, Z => n14883);
   U10164 : BUF_X1 port map( A => n14889, Z => n14884);
   U10165 : BUF_X1 port map( A => n14889, Z => n14885);
   U10166 : BUF_X1 port map( A => n14889, Z => n14886);
   U10167 : BUF_X1 port map( A => n14889, Z => n14887);
   U10168 : BUF_X1 port map( A => n14898, Z => n14891);
   U10169 : BUF_X1 port map( A => n14898, Z => n14892);
   U10170 : BUF_X1 port map( A => n14898, Z => n14893);
   U10171 : BUF_X1 port map( A => n14898, Z => n14894);
   U10172 : BUF_X1 port map( A => n14898, Z => n14895);
   U10173 : BUF_X1 port map( A => n14898, Z => n14896);
   U10174 : BUF_X1 port map( A => n14907, Z => n14900);
   U10175 : BUF_X1 port map( A => n14907, Z => n14901);
   U10176 : BUF_X1 port map( A => n14907, Z => n14902);
   U10177 : BUF_X1 port map( A => n14907, Z => n14903);
   U10178 : BUF_X1 port map( A => n14907, Z => n14904);
   U10179 : BUF_X1 port map( A => n14907, Z => n14905);
   U10180 : BUF_X1 port map( A => n14916, Z => n14909);
   U10181 : BUF_X1 port map( A => n14916, Z => n14910);
   U10182 : BUF_X1 port map( A => n14916, Z => n14911);
   U10183 : BUF_X1 port map( A => n14916, Z => n14912);
   U10184 : BUF_X1 port map( A => n14916, Z => n14913);
   U10185 : BUF_X1 port map( A => n14916, Z => n14914);
   U10186 : BUF_X1 port map( A => n14934, Z => n14927);
   U10187 : BUF_X1 port map( A => n14934, Z => n14928);
   U10188 : BUF_X1 port map( A => n14934, Z => n14929);
   U10189 : BUF_X1 port map( A => n14934, Z => n14930);
   U10190 : BUF_X1 port map( A => n14934, Z => n14931);
   U10191 : BUF_X1 port map( A => n14934, Z => n14932);
   U10192 : BUF_X1 port map( A => n14943, Z => n14936);
   U10193 : BUF_X1 port map( A => n14943, Z => n14937);
   U10194 : BUF_X1 port map( A => n14943, Z => n14938);
   U10195 : BUF_X1 port map( A => n14943, Z => n14939);
   U10196 : BUF_X1 port map( A => n14943, Z => n14940);
   U10197 : BUF_X1 port map( A => n14943, Z => n14941);
   U10198 : BUF_X1 port map( A => n14952, Z => n14945);
   U10199 : BUF_X1 port map( A => n14952, Z => n14946);
   U10200 : BUF_X1 port map( A => n14952, Z => n14947);
   U10201 : BUF_X1 port map( A => n14952, Z => n14948);
   U10202 : BUF_X1 port map( A => n14952, Z => n14949);
   U10203 : BUF_X1 port map( A => n14952, Z => n14950);
   U10204 : BUF_X1 port map( A => n14961, Z => n14954);
   U10205 : BUF_X1 port map( A => n14961, Z => n14955);
   U10206 : BUF_X1 port map( A => n14961, Z => n14956);
   U10207 : BUF_X1 port map( A => n14961, Z => n14957);
   U10208 : BUF_X1 port map( A => n14961, Z => n14958);
   U10209 : BUF_X1 port map( A => n14961, Z => n14959);
   U10210 : BUF_X1 port map( A => n14970, Z => n14963);
   U10211 : BUF_X1 port map( A => n14970, Z => n14964);
   U10212 : BUF_X1 port map( A => n14970, Z => n14965);
   U10213 : BUF_X1 port map( A => n14970, Z => n14966);
   U10214 : BUF_X1 port map( A => n14970, Z => n14967);
   U10215 : BUF_X1 port map( A => n14970, Z => n14968);
   U10216 : BUF_X1 port map( A => n14979, Z => n14972);
   U10217 : BUF_X1 port map( A => n14979, Z => n14973);
   U10218 : BUF_X1 port map( A => n14979, Z => n14974);
   U10219 : BUF_X1 port map( A => n14979, Z => n14975);
   U10220 : BUF_X1 port map( A => n14979, Z => n14976);
   U10221 : BUF_X1 port map( A => n14979, Z => n14977);
   U10222 : BUF_X1 port map( A => n14988, Z => n14981);
   U10223 : BUF_X1 port map( A => n14988, Z => n14982);
   U10224 : BUF_X1 port map( A => n14988, Z => n14983);
   U10225 : BUF_X1 port map( A => n14988, Z => n14984);
   U10226 : BUF_X1 port map( A => n14988, Z => n14985);
   U10227 : BUF_X1 port map( A => n14988, Z => n14986);
   U10228 : BUF_X1 port map( A => n14997, Z => n14990);
   U10229 : BUF_X1 port map( A => n14997, Z => n14991);
   U10230 : BUF_X1 port map( A => n14997, Z => n14992);
   U10231 : BUF_X1 port map( A => n14997, Z => n14993);
   U10232 : BUF_X1 port map( A => n14997, Z => n14994);
   U10233 : BUF_X1 port map( A => n14997, Z => n14995);
   U10234 : BUF_X1 port map( A => n15006, Z => n14999);
   U10235 : BUF_X1 port map( A => n15006, Z => n15000);
   U10236 : BUF_X1 port map( A => n15006, Z => n15001);
   U10237 : BUF_X1 port map( A => n15006, Z => n15002);
   U10238 : BUF_X1 port map( A => n15006, Z => n15003);
   U10239 : BUF_X1 port map( A => n15006, Z => n15004);
   U10240 : BUF_X1 port map( A => n15015, Z => n15008);
   U10241 : BUF_X1 port map( A => n15015, Z => n15009);
   U10242 : BUF_X1 port map( A => n15015, Z => n15010);
   U10243 : BUF_X1 port map( A => n15015, Z => n15011);
   U10244 : BUF_X1 port map( A => n15015, Z => n15012);
   U10245 : BUF_X1 port map( A => n15015, Z => n15013);
   U10246 : BUF_X1 port map( A => n15024, Z => n15017);
   U10247 : BUF_X1 port map( A => n15024, Z => n15018);
   U10248 : BUF_X1 port map( A => n15024, Z => n15019);
   U10249 : BUF_X1 port map( A => n15024, Z => n15020);
   U10250 : BUF_X1 port map( A => n15024, Z => n15021);
   U10251 : BUF_X1 port map( A => n15024, Z => n15022);
   U10252 : BUF_X1 port map( A => n15033, Z => n15026);
   U10253 : BUF_X1 port map( A => n15033, Z => n15027);
   U10254 : BUF_X1 port map( A => n15033, Z => n15028);
   U10255 : BUF_X1 port map( A => n15033, Z => n15029);
   U10256 : BUF_X1 port map( A => n15033, Z => n15030);
   U10257 : BUF_X1 port map( A => n15033, Z => n15031);
   U10258 : BUF_X1 port map( A => n15042, Z => n15035);
   U10259 : BUF_X1 port map( A => n15042, Z => n15036);
   U10260 : BUF_X1 port map( A => n15042, Z => n15037);
   U10261 : BUF_X1 port map( A => n15042, Z => n15038);
   U10262 : BUF_X1 port map( A => n15042, Z => n15039);
   U10263 : BUF_X1 port map( A => n15042, Z => n15040);
   U10264 : BUF_X1 port map( A => n15051, Z => n15044);
   U10265 : BUF_X1 port map( A => n15051, Z => n15045);
   U10266 : BUF_X1 port map( A => n15051, Z => n15046);
   U10267 : BUF_X1 port map( A => n15051, Z => n15047);
   U10268 : BUF_X1 port map( A => n15051, Z => n15048);
   U10269 : BUF_X1 port map( A => n15051, Z => n15049);
   U10270 : BUF_X1 port map( A => n15060, Z => n15053);
   U10271 : BUF_X1 port map( A => n15060, Z => n15054);
   U10272 : BUF_X1 port map( A => n15060, Z => n15055);
   U10273 : BUF_X1 port map( A => n15060, Z => n15056);
   U10274 : BUF_X1 port map( A => n15060, Z => n15057);
   U10275 : BUF_X1 port map( A => n15060, Z => n15058);
   U10276 : BUF_X1 port map( A => n14799, Z => n14798);
   U10277 : BUF_X1 port map( A => n14808, Z => n14807);
   U10278 : BUF_X1 port map( A => n14817, Z => n14816);
   U10279 : BUF_X1 port map( A => n14826, Z => n14825);
   U10280 : BUF_X1 port map( A => n14835, Z => n14834);
   U10281 : BUF_X1 port map( A => n14844, Z => n14843);
   U10282 : BUF_X1 port map( A => n14853, Z => n14852);
   U10283 : BUF_X1 port map( A => n14862, Z => n14861);
   U10284 : BUF_X1 port map( A => n14871, Z => n14870);
   U10285 : BUF_X1 port map( A => n14880, Z => n14879);
   U10286 : BUF_X1 port map( A => n14889, Z => n14888);
   U10287 : BUF_X1 port map( A => n14898, Z => n14897);
   U10288 : BUF_X1 port map( A => n14907, Z => n14906);
   U10289 : BUF_X1 port map( A => n14916, Z => n14915);
   U10290 : BUF_X1 port map( A => n14934, Z => n14933);
   U10291 : BUF_X1 port map( A => n14943, Z => n14942);
   U10292 : BUF_X1 port map( A => n14952, Z => n14951);
   U10293 : BUF_X1 port map( A => n14961, Z => n14960);
   U10294 : BUF_X1 port map( A => n14970, Z => n14969);
   U10295 : BUF_X1 port map( A => n14979, Z => n14978);
   U10296 : BUF_X1 port map( A => n14988, Z => n14987);
   U10297 : BUF_X1 port map( A => n14997, Z => n14996);
   U10298 : BUF_X1 port map( A => n15006, Z => n15005);
   U10299 : BUF_X1 port map( A => n15015, Z => n15014);
   U10300 : BUF_X1 port map( A => n15024, Z => n15023);
   U10301 : BUF_X1 port map( A => n15033, Z => n15032);
   U10302 : BUF_X1 port map( A => n15042, Z => n15041);
   U10303 : BUF_X1 port map( A => n15051, Z => n15050);
   U10304 : BUF_X1 port map( A => n15060, Z => n15059);
   U10305 : AND2_X1 port map( A1 => n14658, A2 => n13182, ZN => n12653);
   U10306 : AND2_X1 port map( A1 => n14756, A2 => n12601, ZN => n12072);
   U10307 : AND2_X1 port map( A1 => n14655, A2 => n13182, ZN => n12656);
   U10308 : AND2_X1 port map( A1 => n14753, A2 => n12601, ZN => n12075);
   U10309 : AND2_X1 port map( A1 => n14044, A2 => n13182, ZN => n12640);
   U10310 : AND2_X1 port map( A1 => n14045, A2 => n12601, ZN => n12059);
   U10311 : INV_X1 port map( A => n11949, ZN => n15162);
   U10312 : OAI21_X1 port map( B1 => n11981, B2 => n11982, A => n15168, ZN => 
                           n11949);
   U10313 : INV_X1 port map( A => n12005, ZN => n14925);
   U10314 : OAI21_X1 port map( B1 => n11982, B2 => n12006, A => n15169, ZN => 
                           n12005);
   U10315 : INV_X1 port map( A => n14780, ZN => n14790);
   U10316 : NOR4_X1 port map( A1 => n13172, A2 => n13173, A3 => n13174, A4 => 
                           n13175, ZN => n13171);
   U10317 : OAI222_X1 port map( A1 => n14094, A2 => n14641, B1 => n13728, B2 =>
                           n14638, C1 => n13832, C2 => n14635, ZN => n13173);
   U10318 : OAI222_X1 port map( A1 => n14118, A2 => n14650, B1 => n13740, B2 =>
                           n14647, C1 => n13844, C2 => n14644, ZN => n13174);
   U10319 : OAI221_X1 port map( B1 => n13812, B2 => n14632, C1 => n14142, C2 =>
                           n14629, A => n13184, ZN => n13172);
   U10320 : NOR4_X1 port map( A1 => n13155, A2 => n13156, A3 => n13157, A4 => 
                           n13158, ZN => n13154);
   U10321 : OAI222_X1 port map( A1 => n14095, A2 => n14641, B1 => n13729, B2 =>
                           n14638, C1 => n13833, C2 => n14635, ZN => n13156);
   U10322 : OAI222_X1 port map( A1 => n14119, A2 => n14650, B1 => n13741, B2 =>
                           n14647, C1 => n13845, C2 => n14644, ZN => n13157);
   U10323 : OAI221_X1 port map( B1 => n13813, B2 => n14632, C1 => n14143, C2 =>
                           n14629, A => n13164, ZN => n13155);
   U10324 : NOR4_X1 port map( A1 => n13138, A2 => n13139, A3 => n13140, A4 => 
                           n13141, ZN => n13137);
   U10325 : OAI222_X1 port map( A1 => n14096, A2 => n14641, B1 => n13730, B2 =>
                           n14638, C1 => n13834, C2 => n14635, ZN => n13139);
   U10326 : OAI222_X1 port map( A1 => n14120, A2 => n14650, B1 => n13742, B2 =>
                           n14647, C1 => n13846, C2 => n14644, ZN => n13140);
   U10327 : OAI221_X1 port map( B1 => n13814, B2 => n14632, C1 => n14144, C2 =>
                           n14629, A => n13147, ZN => n13138);
   U10328 : NOR4_X1 port map( A1 => n13121, A2 => n13122, A3 => n13123, A4 => 
                           n13124, ZN => n13120);
   U10329 : OAI222_X1 port map( A1 => n14097, A2 => n14641, B1 => n13731, B2 =>
                           n14638, C1 => n13835, C2 => n14635, ZN => n13122);
   U10330 : OAI222_X1 port map( A1 => n14121, A2 => n14650, B1 => n13743, B2 =>
                           n14647, C1 => n13847, C2 => n14644, ZN => n13123);
   U10331 : OAI221_X1 port map( B1 => n13815, B2 => n14632, C1 => n14145, C2 =>
                           n14629, A => n13130, ZN => n13121);
   U10332 : NOR4_X1 port map( A1 => n13104, A2 => n13105, A3 => n13106, A4 => 
                           n13107, ZN => n13103);
   U10333 : OAI222_X1 port map( A1 => n14098, A2 => n14641, B1 => n13732, B2 =>
                           n14638, C1 => n13836, C2 => n14635, ZN => n13105);
   U10334 : OAI222_X1 port map( A1 => n14122, A2 => n14650, B1 => n13744, B2 =>
                           n14647, C1 => n13848, C2 => n14644, ZN => n13106);
   U10335 : OAI221_X1 port map( B1 => n13816, B2 => n14632, C1 => n14146, C2 =>
                           n14629, A => n13113, ZN => n13104);
   U10336 : NOR4_X1 port map( A1 => n13087, A2 => n13088, A3 => n13089, A4 => 
                           n13090, ZN => n13086);
   U10337 : OAI222_X1 port map( A1 => n14099, A2 => n14641, B1 => n13733, B2 =>
                           n14638, C1 => n13837, C2 => n14635, ZN => n13088);
   U10338 : OAI222_X1 port map( A1 => n14123, A2 => n14650, B1 => n13745, B2 =>
                           n14647, C1 => n13849, C2 => n14644, ZN => n13089);
   U10339 : OAI221_X1 port map( B1 => n13817, B2 => n14632, C1 => n14147, C2 =>
                           n14629, A => n13096, ZN => n13087);
   U10340 : NOR4_X1 port map( A1 => n13070, A2 => n13071, A3 => n13072, A4 => 
                           n13073, ZN => n13069);
   U10341 : OAI222_X1 port map( A1 => n14100, A2 => n14641, B1 => n13734, B2 =>
                           n14638, C1 => n13838, C2 => n14635, ZN => n13071);
   U10342 : OAI222_X1 port map( A1 => n14124, A2 => n14650, B1 => n13746, B2 =>
                           n14647, C1 => n13850, C2 => n14644, ZN => n13072);
   U10343 : OAI221_X1 port map( B1 => n13818, B2 => n14632, C1 => n14148, C2 =>
                           n14629, A => n13079, ZN => n13070);
   U10344 : NOR4_X1 port map( A1 => n13053, A2 => n13054, A3 => n13055, A4 => 
                           n13056, ZN => n13052);
   U10345 : OAI222_X1 port map( A1 => n14101, A2 => n14641, B1 => n13735, B2 =>
                           n14638, C1 => n13839, C2 => n14635, ZN => n13054);
   U10346 : OAI222_X1 port map( A1 => n14125, A2 => n14650, B1 => n13747, B2 =>
                           n14647, C1 => n13851, C2 => n14644, ZN => n13055);
   U10347 : OAI221_X1 port map( B1 => n13819, B2 => n14632, C1 => n14149, C2 =>
                           n14629, A => n13062, ZN => n13053);
   U10348 : NOR4_X1 port map( A1 => n13036, A2 => n13037, A3 => n13038, A4 => 
                           n13039, ZN => n13035);
   U10349 : OAI222_X1 port map( A1 => n14102, A2 => n14641, B1 => n13736, B2 =>
                           n14638, C1 => n13840, C2 => n14635, ZN => n13037);
   U10350 : OAI222_X1 port map( A1 => n14126, A2 => n14650, B1 => n13748, B2 =>
                           n14647, C1 => n13852, C2 => n14644, ZN => n13038);
   U10351 : OAI221_X1 port map( B1 => n13820, B2 => n14632, C1 => n14150, C2 =>
                           n14629, A => n13045, ZN => n13036);
   U10352 : NOR4_X1 port map( A1 => n13019, A2 => n13020, A3 => n13021, A4 => 
                           n13022, ZN => n13018);
   U10353 : OAI222_X1 port map( A1 => n14103, A2 => n14641, B1 => n13737, B2 =>
                           n14638, C1 => n13841, C2 => n14635, ZN => n13020);
   U10354 : OAI222_X1 port map( A1 => n14127, A2 => n14650, B1 => n13749, B2 =>
                           n14647, C1 => n13853, C2 => n14644, ZN => n13021);
   U10355 : OAI221_X1 port map( B1 => n13821, B2 => n14632, C1 => n14151, C2 =>
                           n14629, A => n13028, ZN => n13019);
   U10356 : NOR4_X1 port map( A1 => n13002, A2 => n13003, A3 => n13004, A4 => 
                           n13005, ZN => n13001);
   U10357 : OAI222_X1 port map( A1 => n14104, A2 => n14641, B1 => n13738, B2 =>
                           n14638, C1 => n13842, C2 => n14635, ZN => n13003);
   U10358 : OAI222_X1 port map( A1 => n14128, A2 => n14650, B1 => n13750, B2 =>
                           n14647, C1 => n13854, C2 => n14644, ZN => n13004);
   U10359 : OAI221_X1 port map( B1 => n13822, B2 => n14632, C1 => n14152, C2 =>
                           n14629, A => n13011, ZN => n13002);
   U10360 : NOR4_X1 port map( A1 => n12985, A2 => n12986, A3 => n12987, A4 => 
                           n12988, ZN => n12984);
   U10361 : OAI222_X1 port map( A1 => n14105, A2 => n14641, B1 => n13739, B2 =>
                           n14638, C1 => n13843, C2 => n14635, ZN => n12986);
   U10362 : OAI222_X1 port map( A1 => n14129, A2 => n14650, B1 => n13751, B2 =>
                           n14647, C1 => n13855, C2 => n14644, ZN => n12987);
   U10363 : OAI221_X1 port map( B1 => n13823, B2 => n14632, C1 => n14153, C2 =>
                           n14629, A => n12994, ZN => n12985);
   U10364 : NOR4_X1 port map( A1 => n12968, A2 => n12969, A3 => n12970, A4 => 
                           n12971, ZN => n12967);
   U10365 : OAI222_X1 port map( A1 => n14106, A2 => n14642, B1 => n13660, B2 =>
                           n14639, C1 => n13768, C2 => n14636, ZN => n12969);
   U10366 : OAI222_X1 port map( A1 => n14130, A2 => n14651, B1 => n13672, B2 =>
                           n14648, C1 => n13780, C2 => n14645, ZN => n12970);
   U10367 : OAI221_X1 port map( B1 => n13712, B2 => n14633, C1 => n14154, C2 =>
                           n14630, A => n12977, ZN => n12968);
   U10368 : NOR4_X1 port map( A1 => n12951, A2 => n12952, A3 => n12953, A4 => 
                           n12954, ZN => n12950);
   U10369 : OAI222_X1 port map( A1 => n14107, A2 => n14642, B1 => n13661, B2 =>
                           n14639, C1 => n13769, C2 => n14636, ZN => n12952);
   U10370 : OAI222_X1 port map( A1 => n14131, A2 => n14651, B1 => n13673, B2 =>
                           n14648, C1 => n13781, C2 => n14645, ZN => n12953);
   U10371 : OAI221_X1 port map( B1 => n13713, B2 => n14633, C1 => n14155, C2 =>
                           n14630, A => n12960, ZN => n12951);
   U10372 : NOR4_X1 port map( A1 => n12934, A2 => n12935, A3 => n12936, A4 => 
                           n12937, ZN => n12933);
   U10373 : OAI222_X1 port map( A1 => n14108, A2 => n14642, B1 => n13662, B2 =>
                           n14639, C1 => n13770, C2 => n14636, ZN => n12935);
   U10374 : OAI222_X1 port map( A1 => n14132, A2 => n14651, B1 => n13674, B2 =>
                           n14648, C1 => n13782, C2 => n14645, ZN => n12936);
   U10375 : OAI221_X1 port map( B1 => n13714, B2 => n14633, C1 => n14156, C2 =>
                           n14630, A => n12943, ZN => n12934);
   U10376 : NOR4_X1 port map( A1 => n12917, A2 => n12918, A3 => n12919, A4 => 
                           n12920, ZN => n12916);
   U10377 : OAI222_X1 port map( A1 => n14109, A2 => n14642, B1 => n13663, B2 =>
                           n14639, C1 => n13771, C2 => n14636, ZN => n12918);
   U10378 : OAI222_X1 port map( A1 => n14133, A2 => n14651, B1 => n13675, B2 =>
                           n14648, C1 => n13783, C2 => n14645, ZN => n12919);
   U10379 : OAI221_X1 port map( B1 => n13715, B2 => n14633, C1 => n14157, C2 =>
                           n14630, A => n12926, ZN => n12917);
   U10380 : NOR4_X1 port map( A1 => n12900, A2 => n12901, A3 => n12902, A4 => 
                           n12903, ZN => n12899);
   U10381 : OAI222_X1 port map( A1 => n14110, A2 => n14642, B1 => n13664, B2 =>
                           n14639, C1 => n13772, C2 => n14636, ZN => n12901);
   U10382 : OAI222_X1 port map( A1 => n14134, A2 => n14651, B1 => n13676, B2 =>
                           n14648, C1 => n13784, C2 => n14645, ZN => n12902);
   U10383 : OAI221_X1 port map( B1 => n13716, B2 => n14633, C1 => n14158, C2 =>
                           n14630, A => n12909, ZN => n12900);
   U10384 : NOR4_X1 port map( A1 => n12883, A2 => n12884, A3 => n12885, A4 => 
                           n12886, ZN => n12882);
   U10385 : OAI222_X1 port map( A1 => n14111, A2 => n14642, B1 => n13665, B2 =>
                           n14639, C1 => n13773, C2 => n14636, ZN => n12884);
   U10386 : OAI222_X1 port map( A1 => n14135, A2 => n14651, B1 => n13677, B2 =>
                           n14648, C1 => n13785, C2 => n14645, ZN => n12885);
   U10387 : OAI221_X1 port map( B1 => n13717, B2 => n14633, C1 => n14159, C2 =>
                           n14630, A => n12892, ZN => n12883);
   U10388 : NOR4_X1 port map( A1 => n12866, A2 => n12867, A3 => n12868, A4 => 
                           n12869, ZN => n12865);
   U10389 : OAI222_X1 port map( A1 => n14112, A2 => n14642, B1 => n13666, B2 =>
                           n14639, C1 => n13774, C2 => n14636, ZN => n12867);
   U10390 : OAI222_X1 port map( A1 => n14136, A2 => n14651, B1 => n13678, B2 =>
                           n14648, C1 => n13786, C2 => n14645, ZN => n12868);
   U10391 : OAI221_X1 port map( B1 => n13718, B2 => n14633, C1 => n14160, C2 =>
                           n14630, A => n12875, ZN => n12866);
   U10392 : NOR4_X1 port map( A1 => n12849, A2 => n12850, A3 => n12851, A4 => 
                           n12852, ZN => n12848);
   U10393 : OAI222_X1 port map( A1 => n14113, A2 => n14642, B1 => n13667, B2 =>
                           n14639, C1 => n13775, C2 => n14636, ZN => n12850);
   U10394 : OAI222_X1 port map( A1 => n14137, A2 => n14651, B1 => n13679, B2 =>
                           n14648, C1 => n13787, C2 => n14645, ZN => n12851);
   U10395 : OAI221_X1 port map( B1 => n13719, B2 => n14633, C1 => n14161, C2 =>
                           n14630, A => n12858, ZN => n12849);
   U10396 : NOR4_X1 port map( A1 => n12832, A2 => n12833, A3 => n12834, A4 => 
                           n12835, ZN => n12831);
   U10397 : OAI222_X1 port map( A1 => n14114, A2 => n14642, B1 => n13668, B2 =>
                           n14639, C1 => n13776, C2 => n14636, ZN => n12833);
   U10398 : OAI222_X1 port map( A1 => n14138, A2 => n14651, B1 => n13680, B2 =>
                           n14648, C1 => n13788, C2 => n14645, ZN => n12834);
   U10399 : OAI221_X1 port map( B1 => n13720, B2 => n14633, C1 => n14162, C2 =>
                           n14630, A => n12841, ZN => n12832);
   U10400 : NOR4_X1 port map( A1 => n12815, A2 => n12816, A3 => n12817, A4 => 
                           n12818, ZN => n12814);
   U10401 : OAI222_X1 port map( A1 => n14115, A2 => n14642, B1 => n13669, B2 =>
                           n14639, C1 => n13777, C2 => n14636, ZN => n12816);
   U10402 : OAI222_X1 port map( A1 => n14139, A2 => n14651, B1 => n13681, B2 =>
                           n14648, C1 => n13789, C2 => n14645, ZN => n12817);
   U10403 : OAI221_X1 port map( B1 => n13721, B2 => n14633, C1 => n14163, C2 =>
                           n14630, A => n12824, ZN => n12815);
   U10404 : NOR4_X1 port map( A1 => n12798, A2 => n12799, A3 => n12800, A4 => 
                           n12801, ZN => n12797);
   U10405 : OAI222_X1 port map( A1 => n14116, A2 => n14642, B1 => n13670, B2 =>
                           n14639, C1 => n13778, C2 => n14636, ZN => n12799);
   U10406 : OAI222_X1 port map( A1 => n14140, A2 => n14651, B1 => n13682, B2 =>
                           n14648, C1 => n13790, C2 => n14645, ZN => n12800);
   U10407 : OAI221_X1 port map( B1 => n13722, B2 => n14633, C1 => n14164, C2 =>
                           n14630, A => n12807, ZN => n12798);
   U10408 : NOR4_X1 port map( A1 => n12781, A2 => n12782, A3 => n12783, A4 => 
                           n12784, ZN => n12780);
   U10409 : OAI222_X1 port map( A1 => n14117, A2 => n14642, B1 => n13671, B2 =>
                           n14639, C1 => n13779, C2 => n14636, ZN => n12782);
   U10410 : OAI222_X1 port map( A1 => n14141, A2 => n14651, B1 => n13683, B2 =>
                           n14648, C1 => n13791, C2 => n14645, ZN => n12783);
   U10411 : OAI221_X1 port map( B1 => n13723, B2 => n14633, C1 => n14165, C2 =>
                           n14630, A => n12790, ZN => n12781);
   U10412 : NOR4_X1 port map( A1 => n12591, A2 => n12592, A3 => n12593, A4 => 
                           n12594, ZN => n12590);
   U10413 : OAI222_X1 port map( A1 => n14094, A2 => n14739, B1 => n13728, B2 =>
                           n14736, C1 => n13832, C2 => n14733, ZN => n12592);
   U10414 : OAI222_X1 port map( A1 => n14118, A2 => n14748, B1 => n13740, B2 =>
                           n14745, C1 => n13844, C2 => n14742, ZN => n12593);
   U10415 : OAI221_X1 port map( B1 => n13812, B2 => n14730, C1 => n14142, C2 =>
                           n14727, A => n12603, ZN => n12591);
   U10416 : NOR4_X1 port map( A1 => n12574, A2 => n12575, A3 => n12576, A4 => 
                           n12577, ZN => n12573);
   U10417 : OAI222_X1 port map( A1 => n14095, A2 => n14739, B1 => n13729, B2 =>
                           n14736, C1 => n13833, C2 => n14733, ZN => n12575);
   U10418 : OAI222_X1 port map( A1 => n14119, A2 => n14748, B1 => n13741, B2 =>
                           n14745, C1 => n13845, C2 => n14742, ZN => n12576);
   U10419 : OAI221_X1 port map( B1 => n13813, B2 => n14730, C1 => n14143, C2 =>
                           n14727, A => n12583, ZN => n12574);
   U10420 : NOR4_X1 port map( A1 => n12557, A2 => n12558, A3 => n12559, A4 => 
                           n12560, ZN => n12556);
   U10421 : OAI222_X1 port map( A1 => n14096, A2 => n14739, B1 => n13730, B2 =>
                           n14736, C1 => n13834, C2 => n14733, ZN => n12558);
   U10422 : OAI222_X1 port map( A1 => n14120, A2 => n14748, B1 => n13742, B2 =>
                           n14745, C1 => n13846, C2 => n14742, ZN => n12559);
   U10423 : OAI221_X1 port map( B1 => n13814, B2 => n14730, C1 => n14144, C2 =>
                           n14727, A => n12566, ZN => n12557);
   U10424 : NOR4_X1 port map( A1 => n12540, A2 => n12541, A3 => n12542, A4 => 
                           n12543, ZN => n12539);
   U10425 : OAI222_X1 port map( A1 => n14097, A2 => n14739, B1 => n13731, B2 =>
                           n14736, C1 => n13835, C2 => n14733, ZN => n12541);
   U10426 : OAI222_X1 port map( A1 => n14121, A2 => n14748, B1 => n13743, B2 =>
                           n14745, C1 => n13847, C2 => n14742, ZN => n12542);
   U10427 : OAI221_X1 port map( B1 => n13815, B2 => n14730, C1 => n14145, C2 =>
                           n14727, A => n12549, ZN => n12540);
   U10428 : NOR4_X1 port map( A1 => n12523, A2 => n12524, A3 => n12525, A4 => 
                           n12526, ZN => n12522);
   U10429 : OAI222_X1 port map( A1 => n14098, A2 => n14739, B1 => n13732, B2 =>
                           n14736, C1 => n13836, C2 => n14733, ZN => n12524);
   U10430 : OAI222_X1 port map( A1 => n14122, A2 => n14748, B1 => n13744, B2 =>
                           n14745, C1 => n13848, C2 => n14742, ZN => n12525);
   U10431 : OAI221_X1 port map( B1 => n13816, B2 => n14730, C1 => n14146, C2 =>
                           n14727, A => n12532, ZN => n12523);
   U10432 : NOR4_X1 port map( A1 => n12506, A2 => n12507, A3 => n12508, A4 => 
                           n12509, ZN => n12505);
   U10433 : OAI222_X1 port map( A1 => n14099, A2 => n14739, B1 => n13733, B2 =>
                           n14736, C1 => n13837, C2 => n14733, ZN => n12507);
   U10434 : OAI222_X1 port map( A1 => n14123, A2 => n14748, B1 => n13745, B2 =>
                           n14745, C1 => n13849, C2 => n14742, ZN => n12508);
   U10435 : OAI221_X1 port map( B1 => n13817, B2 => n14730, C1 => n14147, C2 =>
                           n14727, A => n12515, ZN => n12506);
   U10436 : NOR4_X1 port map( A1 => n12489, A2 => n12490, A3 => n12491, A4 => 
                           n12492, ZN => n12488);
   U10437 : OAI222_X1 port map( A1 => n14100, A2 => n14739, B1 => n13734, B2 =>
                           n14736, C1 => n13838, C2 => n14733, ZN => n12490);
   U10438 : OAI222_X1 port map( A1 => n14124, A2 => n14748, B1 => n13746, B2 =>
                           n14745, C1 => n13850, C2 => n14742, ZN => n12491);
   U10439 : OAI221_X1 port map( B1 => n13818, B2 => n14730, C1 => n14148, C2 =>
                           n14727, A => n12498, ZN => n12489);
   U10440 : NOR4_X1 port map( A1 => n12472, A2 => n12473, A3 => n12474, A4 => 
                           n12475, ZN => n12471);
   U10441 : OAI222_X1 port map( A1 => n14101, A2 => n14739, B1 => n13735, B2 =>
                           n14736, C1 => n13839, C2 => n14733, ZN => n12473);
   U10442 : OAI222_X1 port map( A1 => n14125, A2 => n14748, B1 => n13747, B2 =>
                           n14745, C1 => n13851, C2 => n14742, ZN => n12474);
   U10443 : OAI221_X1 port map( B1 => n13819, B2 => n14730, C1 => n14149, C2 =>
                           n14727, A => n12481, ZN => n12472);
   U10444 : NOR4_X1 port map( A1 => n12455, A2 => n12456, A3 => n12457, A4 => 
                           n12458, ZN => n12454);
   U10445 : OAI222_X1 port map( A1 => n14102, A2 => n14739, B1 => n13736, B2 =>
                           n14736, C1 => n13840, C2 => n14733, ZN => n12456);
   U10446 : OAI222_X1 port map( A1 => n14126, A2 => n14748, B1 => n13748, B2 =>
                           n14745, C1 => n13852, C2 => n14742, ZN => n12457);
   U10447 : OAI221_X1 port map( B1 => n13820, B2 => n14730, C1 => n14150, C2 =>
                           n14727, A => n12464, ZN => n12455);
   U10448 : NOR4_X1 port map( A1 => n12438, A2 => n12439, A3 => n12440, A4 => 
                           n12441, ZN => n12437);
   U10449 : OAI222_X1 port map( A1 => n14103, A2 => n14739, B1 => n13737, B2 =>
                           n14736, C1 => n13841, C2 => n14733, ZN => n12439);
   U10450 : OAI222_X1 port map( A1 => n14127, A2 => n14748, B1 => n13749, B2 =>
                           n14745, C1 => n13853, C2 => n14742, ZN => n12440);
   U10451 : OAI221_X1 port map( B1 => n13821, B2 => n14730, C1 => n14151, C2 =>
                           n14727, A => n12447, ZN => n12438);
   U10452 : NOR4_X1 port map( A1 => n12421, A2 => n12422, A3 => n12423, A4 => 
                           n12424, ZN => n12420);
   U10453 : OAI222_X1 port map( A1 => n14104, A2 => n14739, B1 => n13738, B2 =>
                           n14736, C1 => n13842, C2 => n14733, ZN => n12422);
   U10454 : OAI222_X1 port map( A1 => n14128, A2 => n14748, B1 => n13750, B2 =>
                           n14745, C1 => n13854, C2 => n14742, ZN => n12423);
   U10455 : OAI221_X1 port map( B1 => n13822, B2 => n14730, C1 => n14152, C2 =>
                           n14727, A => n12430, ZN => n12421);
   U10456 : NOR4_X1 port map( A1 => n12404, A2 => n12405, A3 => n12406, A4 => 
                           n12407, ZN => n12403);
   U10457 : OAI222_X1 port map( A1 => n14105, A2 => n14739, B1 => n13739, B2 =>
                           n14736, C1 => n13843, C2 => n14733, ZN => n12405);
   U10458 : OAI222_X1 port map( A1 => n14129, A2 => n14748, B1 => n13751, B2 =>
                           n14745, C1 => n13855, C2 => n14742, ZN => n12406);
   U10459 : OAI221_X1 port map( B1 => n13823, B2 => n14730, C1 => n14153, C2 =>
                           n14727, A => n12413, ZN => n12404);
   U10460 : NOR4_X1 port map( A1 => n12387, A2 => n12388, A3 => n12389, A4 => 
                           n12390, ZN => n12386);
   U10461 : OAI222_X1 port map( A1 => n14106, A2 => n14740, B1 => n13660, B2 =>
                           n14737, C1 => n13768, C2 => n14734, ZN => n12388);
   U10462 : OAI222_X1 port map( A1 => n14130, A2 => n14749, B1 => n13672, B2 =>
                           n14746, C1 => n13780, C2 => n14743, ZN => n12389);
   U10463 : OAI221_X1 port map( B1 => n13712, B2 => n14731, C1 => n14154, C2 =>
                           n14728, A => n12396, ZN => n12387);
   U10464 : NOR4_X1 port map( A1 => n12370, A2 => n12371, A3 => n12372, A4 => 
                           n12373, ZN => n12369);
   U10465 : OAI222_X1 port map( A1 => n14107, A2 => n14740, B1 => n13661, B2 =>
                           n14737, C1 => n13769, C2 => n14734, ZN => n12371);
   U10466 : OAI222_X1 port map( A1 => n14131, A2 => n14749, B1 => n13673, B2 =>
                           n14746, C1 => n13781, C2 => n14743, ZN => n12372);
   U10467 : OAI221_X1 port map( B1 => n13713, B2 => n14731, C1 => n14155, C2 =>
                           n14728, A => n12379, ZN => n12370);
   U10468 : NOR4_X1 port map( A1 => n12353, A2 => n12354, A3 => n12355, A4 => 
                           n12356, ZN => n12352);
   U10469 : OAI222_X1 port map( A1 => n14108, A2 => n14740, B1 => n13662, B2 =>
                           n14737, C1 => n13770, C2 => n14734, ZN => n12354);
   U10470 : OAI222_X1 port map( A1 => n14132, A2 => n14749, B1 => n13674, B2 =>
                           n14746, C1 => n13782, C2 => n14743, ZN => n12355);
   U10471 : OAI221_X1 port map( B1 => n13714, B2 => n14731, C1 => n14156, C2 =>
                           n14728, A => n12362, ZN => n12353);
   U10472 : NOR4_X1 port map( A1 => n12336, A2 => n12337, A3 => n12338, A4 => 
                           n12339, ZN => n12335);
   U10473 : OAI222_X1 port map( A1 => n14109, A2 => n14740, B1 => n13663, B2 =>
                           n14737, C1 => n13771, C2 => n14734, ZN => n12337);
   U10474 : OAI222_X1 port map( A1 => n14133, A2 => n14749, B1 => n13675, B2 =>
                           n14746, C1 => n13783, C2 => n14743, ZN => n12338);
   U10475 : OAI221_X1 port map( B1 => n13715, B2 => n14731, C1 => n14157, C2 =>
                           n14728, A => n12345, ZN => n12336);
   U10476 : NOR4_X1 port map( A1 => n12319, A2 => n12320, A3 => n12321, A4 => 
                           n12322, ZN => n12318);
   U10477 : OAI222_X1 port map( A1 => n14110, A2 => n14740, B1 => n13664, B2 =>
                           n14737, C1 => n13772, C2 => n14734, ZN => n12320);
   U10478 : OAI222_X1 port map( A1 => n14134, A2 => n14749, B1 => n13676, B2 =>
                           n14746, C1 => n13784, C2 => n14743, ZN => n12321);
   U10479 : OAI221_X1 port map( B1 => n13716, B2 => n14731, C1 => n14158, C2 =>
                           n14728, A => n12328, ZN => n12319);
   U10480 : NOR4_X1 port map( A1 => n12302, A2 => n12303, A3 => n12304, A4 => 
                           n12305, ZN => n12301);
   U10481 : OAI222_X1 port map( A1 => n14111, A2 => n14740, B1 => n13665, B2 =>
                           n14737, C1 => n13773, C2 => n14734, ZN => n12303);
   U10482 : OAI222_X1 port map( A1 => n14135, A2 => n14749, B1 => n13677, B2 =>
                           n14746, C1 => n13785, C2 => n14743, ZN => n12304);
   U10483 : OAI221_X1 port map( B1 => n13717, B2 => n14731, C1 => n14159, C2 =>
                           n14728, A => n12311, ZN => n12302);
   U10484 : NOR4_X1 port map( A1 => n12285, A2 => n12286, A3 => n12287, A4 => 
                           n12288, ZN => n12284);
   U10485 : OAI222_X1 port map( A1 => n14112, A2 => n14740, B1 => n13666, B2 =>
                           n14737, C1 => n13774, C2 => n14734, ZN => n12286);
   U10486 : OAI222_X1 port map( A1 => n14136, A2 => n14749, B1 => n13678, B2 =>
                           n14746, C1 => n13786, C2 => n14743, ZN => n12287);
   U10487 : OAI221_X1 port map( B1 => n13718, B2 => n14731, C1 => n14160, C2 =>
                           n14728, A => n12294, ZN => n12285);
   U10488 : NOR4_X1 port map( A1 => n12268, A2 => n12269, A3 => n12270, A4 => 
                           n12271, ZN => n12267);
   U10489 : OAI222_X1 port map( A1 => n14113, A2 => n14740, B1 => n13667, B2 =>
                           n14737, C1 => n13775, C2 => n14734, ZN => n12269);
   U10490 : OAI222_X1 port map( A1 => n14137, A2 => n14749, B1 => n13679, B2 =>
                           n14746, C1 => n13787, C2 => n14743, ZN => n12270);
   U10491 : OAI221_X1 port map( B1 => n13719, B2 => n14731, C1 => n14161, C2 =>
                           n14728, A => n12277, ZN => n12268);
   U10492 : NOR4_X1 port map( A1 => n12251, A2 => n12252, A3 => n12253, A4 => 
                           n12254, ZN => n12250);
   U10493 : OAI222_X1 port map( A1 => n14114, A2 => n14740, B1 => n13668, B2 =>
                           n14737, C1 => n13776, C2 => n14734, ZN => n12252);
   U10494 : OAI222_X1 port map( A1 => n14138, A2 => n14749, B1 => n13680, B2 =>
                           n14746, C1 => n13788, C2 => n14743, ZN => n12253);
   U10495 : OAI221_X1 port map( B1 => n13720, B2 => n14731, C1 => n14162, C2 =>
                           n14728, A => n12260, ZN => n12251);
   U10496 : NOR4_X1 port map( A1 => n12234, A2 => n12235, A3 => n12236, A4 => 
                           n12237, ZN => n12233);
   U10497 : OAI222_X1 port map( A1 => n14115, A2 => n14740, B1 => n13669, B2 =>
                           n14737, C1 => n13777, C2 => n14734, ZN => n12235);
   U10498 : OAI222_X1 port map( A1 => n14139, A2 => n14749, B1 => n13681, B2 =>
                           n14746, C1 => n13789, C2 => n14743, ZN => n12236);
   U10499 : OAI221_X1 port map( B1 => n13721, B2 => n14731, C1 => n14163, C2 =>
                           n14728, A => n12243, ZN => n12234);
   U10500 : NOR4_X1 port map( A1 => n12217, A2 => n12218, A3 => n12219, A4 => 
                           n12220, ZN => n12216);
   U10501 : OAI222_X1 port map( A1 => n14116, A2 => n14740, B1 => n13670, B2 =>
                           n14737, C1 => n13778, C2 => n14734, ZN => n12218);
   U10502 : OAI222_X1 port map( A1 => n14140, A2 => n14749, B1 => n13682, B2 =>
                           n14746, C1 => n13790, C2 => n14743, ZN => n12219);
   U10503 : OAI221_X1 port map( B1 => n13722, B2 => n14731, C1 => n14164, C2 =>
                           n14728, A => n12226, ZN => n12217);
   U10504 : NOR4_X1 port map( A1 => n12200, A2 => n12201, A3 => n12202, A4 => 
                           n12203, ZN => n12199);
   U10505 : OAI222_X1 port map( A1 => n14117, A2 => n14740, B1 => n13671, B2 =>
                           n14737, C1 => n13779, C2 => n14734, ZN => n12201);
   U10506 : OAI222_X1 port map( A1 => n14141, A2 => n14749, B1 => n13683, B2 =>
                           n14746, C1 => n13791, C2 => n14743, ZN => n12202);
   U10507 : OAI221_X1 port map( B1 => n13723, B2 => n14731, C1 => n14165, C2 =>
                           n14728, A => n12209, ZN => n12200);
   U10508 : NOR4_X1 port map( A1 => n12764, A2 => n12765, A3 => n12766, A4 => 
                           n12767, ZN => n12763);
   U10509 : OAI222_X1 port map( A1 => n13856, A2 => n14643, B1 => n13644, B2 =>
                           n14640, C1 => n13752, C2 => n14637, ZN => n12765);
   U10510 : OAI222_X1 port map( A1 => n13864, A2 => n14652, B1 => n13652, B2 =>
                           n14649, C1 => n13760, C2 => n14646, ZN => n12766);
   U10511 : OAI221_X1 port map( B1 => n13704, B2 => n14634, C1 => n13872, C2 =>
                           n14631, A => n12773, ZN => n12764);
   U10512 : NOR4_X1 port map( A1 => n12747, A2 => n12748, A3 => n12749, A4 => 
                           n12750, ZN => n12746);
   U10513 : OAI222_X1 port map( A1 => n13857, A2 => n14643, B1 => n13645, B2 =>
                           n14640, C1 => n13753, C2 => n14637, ZN => n12748);
   U10514 : OAI222_X1 port map( A1 => n13865, A2 => n14652, B1 => n13653, B2 =>
                           n14649, C1 => n13761, C2 => n14646, ZN => n12749);
   U10515 : OAI221_X1 port map( B1 => n13705, B2 => n14634, C1 => n13873, C2 =>
                           n14631, A => n12756, ZN => n12747);
   U10516 : NOR4_X1 port map( A1 => n12730, A2 => n12731, A3 => n12732, A4 => 
                           n12733, ZN => n12729);
   U10517 : OAI222_X1 port map( A1 => n13858, A2 => n14643, B1 => n13646, B2 =>
                           n14640, C1 => n13754, C2 => n14637, ZN => n12731);
   U10518 : OAI222_X1 port map( A1 => n13866, A2 => n14652, B1 => n13654, B2 =>
                           n14649, C1 => n13762, C2 => n14646, ZN => n12732);
   U10519 : OAI221_X1 port map( B1 => n13706, B2 => n14634, C1 => n13874, C2 =>
                           n14631, A => n12739, ZN => n12730);
   U10520 : NOR4_X1 port map( A1 => n12713, A2 => n12714, A3 => n12715, A4 => 
                           n12716, ZN => n12712);
   U10521 : OAI222_X1 port map( A1 => n13859, A2 => n14643, B1 => n13647, B2 =>
                           n14640, C1 => n13755, C2 => n14637, ZN => n12714);
   U10522 : OAI222_X1 port map( A1 => n13867, A2 => n14652, B1 => n13655, B2 =>
                           n14649, C1 => n13763, C2 => n14646, ZN => n12715);
   U10523 : OAI221_X1 port map( B1 => n13707, B2 => n14634, C1 => n13875, C2 =>
                           n14631, A => n12722, ZN => n12713);
   U10524 : NOR4_X1 port map( A1 => n12696, A2 => n12697, A3 => n12698, A4 => 
                           n12699, ZN => n12695);
   U10525 : OAI222_X1 port map( A1 => n13860, A2 => n14643, B1 => n13648, B2 =>
                           n14640, C1 => n13756, C2 => n14637, ZN => n12697);
   U10526 : OAI222_X1 port map( A1 => n13868, A2 => n14652, B1 => n13656, B2 =>
                           n14649, C1 => n13764, C2 => n14646, ZN => n12698);
   U10527 : OAI221_X1 port map( B1 => n13708, B2 => n14634, C1 => n13876, C2 =>
                           n14631, A => n12705, ZN => n12696);
   U10528 : NOR4_X1 port map( A1 => n12679, A2 => n12680, A3 => n12681, A4 => 
                           n12682, ZN => n12678);
   U10529 : OAI222_X1 port map( A1 => n13861, A2 => n14643, B1 => n13649, B2 =>
                           n14640, C1 => n13757, C2 => n14637, ZN => n12680);
   U10530 : OAI222_X1 port map( A1 => n13869, A2 => n14652, B1 => n13657, B2 =>
                           n14649, C1 => n13765, C2 => n14646, ZN => n12681);
   U10531 : OAI221_X1 port map( B1 => n13709, B2 => n14634, C1 => n13877, C2 =>
                           n14631, A => n12688, ZN => n12679);
   U10532 : NOR4_X1 port map( A1 => n12662, A2 => n12663, A3 => n12664, A4 => 
                           n12665, ZN => n12661);
   U10533 : OAI222_X1 port map( A1 => n13862, A2 => n14643, B1 => n13650, B2 =>
                           n14640, C1 => n13758, C2 => n14637, ZN => n12663);
   U10534 : OAI222_X1 port map( A1 => n13870, A2 => n14652, B1 => n13658, B2 =>
                           n14649, C1 => n13766, C2 => n14646, ZN => n12664);
   U10535 : OAI221_X1 port map( B1 => n13710, B2 => n14634, C1 => n13878, C2 =>
                           n14631, A => n12671, ZN => n12662);
   U10536 : NOR4_X1 port map( A1 => n12611, A2 => n12612, A3 => n12613, A4 => 
                           n12614, ZN => n12610);
   U10537 : OAI222_X1 port map( A1 => n13863, A2 => n14643, B1 => n13651, B2 =>
                           n14640, C1 => n13759, C2 => n14637, ZN => n12612);
   U10538 : OAI222_X1 port map( A1 => n13871, A2 => n14652, B1 => n13659, B2 =>
                           n14649, C1 => n13767, C2 => n14646, ZN => n12613);
   U10539 : OAI221_X1 port map( B1 => n13711, B2 => n14634, C1 => n13879, C2 =>
                           n14631, A => n12639, ZN => n12611);
   U10540 : NOR4_X1 port map( A1 => n12183, A2 => n12184, A3 => n12185, A4 => 
                           n12186, ZN => n12182);
   U10541 : OAI222_X1 port map( A1 => n13856, A2 => n14741, B1 => n13644, B2 =>
                           n14738, C1 => n13752, C2 => n14735, ZN => n12184);
   U10542 : OAI222_X1 port map( A1 => n13864, A2 => n14750, B1 => n13652, B2 =>
                           n14747, C1 => n13760, C2 => n14744, ZN => n12185);
   U10543 : OAI221_X1 port map( B1 => n13704, B2 => n14732, C1 => n13872, C2 =>
                           n14729, A => n12192, ZN => n12183);
   U10544 : NOR4_X1 port map( A1 => n12166, A2 => n12167, A3 => n12168, A4 => 
                           n12169, ZN => n12165);
   U10545 : OAI222_X1 port map( A1 => n13857, A2 => n14741, B1 => n13645, B2 =>
                           n14738, C1 => n13753, C2 => n14735, ZN => n12167);
   U10546 : OAI222_X1 port map( A1 => n13865, A2 => n14750, B1 => n13653, B2 =>
                           n14747, C1 => n13761, C2 => n14744, ZN => n12168);
   U10547 : OAI221_X1 port map( B1 => n13705, B2 => n14732, C1 => n13873, C2 =>
                           n14729, A => n12175, ZN => n12166);
   U10548 : NOR4_X1 port map( A1 => n12149, A2 => n12150, A3 => n12151, A4 => 
                           n12152, ZN => n12148);
   U10549 : OAI222_X1 port map( A1 => n13858, A2 => n14741, B1 => n13646, B2 =>
                           n14738, C1 => n13754, C2 => n14735, ZN => n12150);
   U10550 : OAI222_X1 port map( A1 => n13866, A2 => n14750, B1 => n13654, B2 =>
                           n14747, C1 => n13762, C2 => n14744, ZN => n12151);
   U10551 : OAI221_X1 port map( B1 => n13706, B2 => n14732, C1 => n13874, C2 =>
                           n14729, A => n12158, ZN => n12149);
   U10552 : NOR4_X1 port map( A1 => n12132, A2 => n12133, A3 => n12134, A4 => 
                           n12135, ZN => n12131);
   U10553 : OAI222_X1 port map( A1 => n13859, A2 => n14741, B1 => n13647, B2 =>
                           n14738, C1 => n13755, C2 => n14735, ZN => n12133);
   U10554 : OAI222_X1 port map( A1 => n13867, A2 => n14750, B1 => n13655, B2 =>
                           n14747, C1 => n13763, C2 => n14744, ZN => n12134);
   U10555 : OAI221_X1 port map( B1 => n13707, B2 => n14732, C1 => n13875, C2 =>
                           n14729, A => n12141, ZN => n12132);
   U10556 : NOR4_X1 port map( A1 => n12115, A2 => n12116, A3 => n12117, A4 => 
                           n12118, ZN => n12114);
   U10557 : OAI222_X1 port map( A1 => n13860, A2 => n14741, B1 => n13648, B2 =>
                           n14738, C1 => n13756, C2 => n14735, ZN => n12116);
   U10558 : OAI222_X1 port map( A1 => n13868, A2 => n14750, B1 => n13656, B2 =>
                           n14747, C1 => n13764, C2 => n14744, ZN => n12117);
   U10559 : OAI221_X1 port map( B1 => n13708, B2 => n14732, C1 => n13876, C2 =>
                           n14729, A => n12124, ZN => n12115);
   U10560 : NOR4_X1 port map( A1 => n12098, A2 => n12099, A3 => n12100, A4 => 
                           n12101, ZN => n12097);
   U10561 : OAI222_X1 port map( A1 => n13861, A2 => n14741, B1 => n13649, B2 =>
                           n14738, C1 => n13757, C2 => n14735, ZN => n12099);
   U10562 : OAI222_X1 port map( A1 => n13869, A2 => n14750, B1 => n13657, B2 =>
                           n14747, C1 => n13765, C2 => n14744, ZN => n12100);
   U10563 : OAI221_X1 port map( B1 => n13709, B2 => n14732, C1 => n13877, C2 =>
                           n14729, A => n12107, ZN => n12098);
   U10564 : NOR4_X1 port map( A1 => n12081, A2 => n12082, A3 => n12083, A4 => 
                           n12084, ZN => n12080);
   U10565 : OAI222_X1 port map( A1 => n13862, A2 => n14741, B1 => n13650, B2 =>
                           n14738, C1 => n13758, C2 => n14735, ZN => n12082);
   U10566 : OAI222_X1 port map( A1 => n13870, A2 => n14750, B1 => n13658, B2 =>
                           n14747, C1 => n13766, C2 => n14744, ZN => n12083);
   U10567 : OAI221_X1 port map( B1 => n13710, B2 => n14732, C1 => n13878, C2 =>
                           n14729, A => n12090, ZN => n12081);
   U10568 : NOR4_X1 port map( A1 => n12030, A2 => n12031, A3 => n12032, A4 => 
                           n12033, ZN => n12029);
   U10569 : OAI222_X1 port map( A1 => n13863, A2 => n14741, B1 => n13651, B2 =>
                           n14738, C1 => n13759, C2 => n14735, ZN => n12031);
   U10570 : OAI222_X1 port map( A1 => n13871, A2 => n14750, B1 => n13659, B2 =>
                           n14747, C1 => n13767, C2 => n14744, ZN => n12032);
   U10571 : OAI221_X1 port map( B1 => n13711, B2 => n14732, C1 => n13879, C2 =>
                           n14729, A => n12058, ZN => n12030);
   U10572 : OAI22_X1 port map( A1 => n13684, A2 => n14619, B1 => n13804, B2 => 
                           n14616, ZN => n12775);
   U10573 : OAI22_X1 port map( A1 => n13685, A2 => n14619, B1 => n13805, B2 => 
                           n14616, ZN => n12758);
   U10574 : OAI22_X1 port map( A1 => n13686, A2 => n14619, B1 => n13806, B2 => 
                           n14616, ZN => n12741);
   U10575 : OAI22_X1 port map( A1 => n13687, A2 => n14619, B1 => n13807, B2 => 
                           n14616, ZN => n12724);
   U10576 : OAI22_X1 port map( A1 => n13688, A2 => n14619, B1 => n13808, B2 => 
                           n14616, ZN => n12707);
   U10577 : OAI22_X1 port map( A1 => n13689, A2 => n14619, B1 => n13809, B2 => 
                           n14616, ZN => n12690);
   U10578 : OAI22_X1 port map( A1 => n13690, A2 => n14619, B1 => n13810, B2 => 
                           n14616, ZN => n12673);
   U10579 : OAI22_X1 port map( A1 => n13691, A2 => n14619, B1 => n13811, B2 => 
                           n14616, ZN => n12644);
   U10580 : OAI22_X1 port map( A1 => n13684, A2 => n14717, B1 => n13804, B2 => 
                           n14714, ZN => n12194);
   U10581 : OAI22_X1 port map( A1 => n13685, A2 => n14717, B1 => n13805, B2 => 
                           n14714, ZN => n12177);
   U10582 : OAI22_X1 port map( A1 => n13686, A2 => n14717, B1 => n13806, B2 => 
                           n14714, ZN => n12160);
   U10583 : OAI22_X1 port map( A1 => n13687, A2 => n14717, B1 => n13807, B2 => 
                           n14714, ZN => n12143);
   U10584 : OAI22_X1 port map( A1 => n13688, A2 => n14717, B1 => n13808, B2 => 
                           n14714, ZN => n12126);
   U10585 : OAI22_X1 port map( A1 => n13689, A2 => n14717, B1 => n13809, B2 => 
                           n14714, ZN => n12109);
   U10586 : OAI22_X1 port map( A1 => n13690, A2 => n14717, B1 => n13810, B2 => 
                           n14714, ZN => n12092);
   U10587 : OAI22_X1 port map( A1 => n13691, A2 => n14717, B1 => n13811, B2 => 
                           n14714, ZN => n12063);
   U10588 : OAI22_X1 port map( A1 => n13792, A2 => n14617, B1 => n14046, B2 => 
                           n14614, ZN => n13186);
   U10589 : OAI22_X1 port map( A1 => n13793, A2 => n14617, B1 => n14047, B2 => 
                           n14614, ZN => n13166);
   U10590 : OAI22_X1 port map( A1 => n13794, A2 => n14617, B1 => n14048, B2 => 
                           n14614, ZN => n13149);
   U10591 : OAI22_X1 port map( A1 => n13795, A2 => n14617, B1 => n14049, B2 => 
                           n14614, ZN => n13132);
   U10592 : OAI22_X1 port map( A1 => n13796, A2 => n14617, B1 => n14050, B2 => 
                           n14614, ZN => n13115);
   U10593 : OAI22_X1 port map( A1 => n13797, A2 => n14617, B1 => n14051, B2 => 
                           n14614, ZN => n13098);
   U10594 : OAI22_X1 port map( A1 => n13798, A2 => n14617, B1 => n14052, B2 => 
                           n14614, ZN => n13081);
   U10595 : OAI22_X1 port map( A1 => n13799, A2 => n14617, B1 => n14053, B2 => 
                           n14614, ZN => n13064);
   U10596 : OAI22_X1 port map( A1 => n13800, A2 => n14617, B1 => n14054, B2 => 
                           n14614, ZN => n13047);
   U10597 : OAI22_X1 port map( A1 => n13801, A2 => n14617, B1 => n14055, B2 => 
                           n14614, ZN => n13030);
   U10598 : OAI22_X1 port map( A1 => n13802, A2 => n14617, B1 => n14056, B2 => 
                           n14614, ZN => n13013);
   U10599 : OAI22_X1 port map( A1 => n13803, A2 => n14617, B1 => n14057, B2 => 
                           n14614, ZN => n12996);
   U10600 : OAI22_X1 port map( A1 => n13692, A2 => n14618, B1 => n14058, B2 => 
                           n14615, ZN => n12979);
   U10601 : OAI22_X1 port map( A1 => n13693, A2 => n14618, B1 => n14059, B2 => 
                           n14615, ZN => n12962);
   U10602 : OAI22_X1 port map( A1 => n13694, A2 => n14618, B1 => n14060, B2 => 
                           n14615, ZN => n12945);
   U10603 : OAI22_X1 port map( A1 => n13695, A2 => n14618, B1 => n14061, B2 => 
                           n14615, ZN => n12928);
   U10604 : OAI22_X1 port map( A1 => n13696, A2 => n14618, B1 => n14062, B2 => 
                           n14615, ZN => n12911);
   U10605 : OAI22_X1 port map( A1 => n13697, A2 => n14618, B1 => n14063, B2 => 
                           n14615, ZN => n12894);
   U10606 : OAI22_X1 port map( A1 => n13698, A2 => n14618, B1 => n14064, B2 => 
                           n14615, ZN => n12877);
   U10607 : OAI22_X1 port map( A1 => n13699, A2 => n14618, B1 => n14065, B2 => 
                           n14615, ZN => n12860);
   U10608 : OAI22_X1 port map( A1 => n13700, A2 => n14618, B1 => n14066, B2 => 
                           n14615, ZN => n12843);
   U10609 : OAI22_X1 port map( A1 => n13701, A2 => n14618, B1 => n14067, B2 => 
                           n14615, ZN => n12826);
   U10610 : OAI22_X1 port map( A1 => n13702, A2 => n14618, B1 => n14068, B2 => 
                           n14615, ZN => n12809);
   U10611 : OAI22_X1 port map( A1 => n13703, A2 => n14618, B1 => n14069, B2 => 
                           n14615, ZN => n12792);
   U10612 : OAI22_X1 port map( A1 => n13792, A2 => n14715, B1 => n14046, B2 => 
                           n14712, ZN => n12605);
   U10613 : OAI22_X1 port map( A1 => n13793, A2 => n14715, B1 => n14047, B2 => 
                           n14712, ZN => n12585);
   U10614 : OAI22_X1 port map( A1 => n13794, A2 => n14715, B1 => n14048, B2 => 
                           n14712, ZN => n12568);
   U10615 : OAI22_X1 port map( A1 => n13795, A2 => n14715, B1 => n14049, B2 => 
                           n14712, ZN => n12551);
   U10616 : OAI22_X1 port map( A1 => n13796, A2 => n14715, B1 => n14050, B2 => 
                           n14712, ZN => n12534);
   U10617 : OAI22_X1 port map( A1 => n13797, A2 => n14715, B1 => n14051, B2 => 
                           n14712, ZN => n12517);
   U10618 : OAI22_X1 port map( A1 => n13798, A2 => n14715, B1 => n14052, B2 => 
                           n14712, ZN => n12500);
   U10619 : OAI22_X1 port map( A1 => n13799, A2 => n14715, B1 => n14053, B2 => 
                           n14712, ZN => n12483);
   U10620 : OAI22_X1 port map( A1 => n13800, A2 => n14715, B1 => n14054, B2 => 
                           n14712, ZN => n12466);
   U10621 : OAI22_X1 port map( A1 => n13801, A2 => n14715, B1 => n14055, B2 => 
                           n14712, ZN => n12449);
   U10622 : OAI22_X1 port map( A1 => n13802, A2 => n14715, B1 => n14056, B2 => 
                           n14712, ZN => n12432);
   U10623 : OAI22_X1 port map( A1 => n13803, A2 => n14715, B1 => n14057, B2 => 
                           n14712, ZN => n12415);
   U10624 : OAI22_X1 port map( A1 => n13692, A2 => n14716, B1 => n14058, B2 => 
                           n14713, ZN => n12398);
   U10625 : OAI22_X1 port map( A1 => n13693, A2 => n14716, B1 => n14059, B2 => 
                           n14713, ZN => n12381);
   U10626 : OAI22_X1 port map( A1 => n13694, A2 => n14716, B1 => n14060, B2 => 
                           n14713, ZN => n12364);
   U10627 : OAI22_X1 port map( A1 => n13695, A2 => n14716, B1 => n14061, B2 => 
                           n14713, ZN => n12347);
   U10628 : OAI22_X1 port map( A1 => n13696, A2 => n14716, B1 => n14062, B2 => 
                           n14713, ZN => n12330);
   U10629 : OAI22_X1 port map( A1 => n13697, A2 => n14716, B1 => n14063, B2 => 
                           n14713, ZN => n12313);
   U10630 : OAI22_X1 port map( A1 => n13698, A2 => n14716, B1 => n14064, B2 => 
                           n14713, ZN => n12296);
   U10631 : OAI22_X1 port map( A1 => n13699, A2 => n14716, B1 => n14065, B2 => 
                           n14713, ZN => n12279);
   U10632 : OAI22_X1 port map( A1 => n13700, A2 => n14716, B1 => n14066, B2 => 
                           n14713, ZN => n12262);
   U10633 : OAI22_X1 port map( A1 => n13701, A2 => n14716, B1 => n14067, B2 => 
                           n14713, ZN => n12245);
   U10634 : OAI22_X1 port map( A1 => n13702, A2 => n14716, B1 => n14068, B2 => 
                           n14713, ZN => n12228);
   U10635 : OAI22_X1 port map( A1 => n13703, A2 => n14716, B1 => n14069, B2 => 
                           n14713, ZN => n12211);
   U10636 : OAI22_X1 port map( A1 => n14859, A2 => n15134, B1 => n12015, B2 => 
                           n13892, ZN => n1622);
   U10637 : OAI22_X1 port map( A1 => n14860, A2 => n15137, B1 => n12015, B2 => 
                           n13894, ZN => n1623);
   U10638 : OAI22_X1 port map( A1 => n14860, A2 => n15140, B1 => n12015, B2 => 
                           n13896, ZN => n1624);
   U10639 : OAI22_X1 port map( A1 => n14860, A2 => n15143, B1 => n12015, B2 => 
                           n13898, ZN => n1625);
   U10640 : OAI22_X1 port map( A1 => n14860, A2 => n15146, B1 => n12015, B2 => 
                           n13900, ZN => n1626);
   U10641 : OAI22_X1 port map( A1 => n14860, A2 => n15149, B1 => n12015, B2 => 
                           n13902, ZN => n1627);
   U10642 : OAI22_X1 port map( A1 => n14861, A2 => n15152, B1 => n12015, B2 => 
                           n13904, ZN => n1628);
   U10643 : OAI22_X1 port map( A1 => n14861, A2 => n15164, B1 => n12015, B2 => 
                           n13906, ZN => n1629);
   U10644 : OAI22_X1 port map( A1 => n14868, A2 => n15134, B1 => n12014, B2 => 
                           n13684, ZN => n1654);
   U10645 : OAI22_X1 port map( A1 => n14869, A2 => n15137, B1 => n12014, B2 => 
                           n13685, ZN => n1655);
   U10646 : OAI22_X1 port map( A1 => n14869, A2 => n15140, B1 => n12014, B2 => 
                           n13686, ZN => n1656);
   U10647 : OAI22_X1 port map( A1 => n14869, A2 => n15143, B1 => n12014, B2 => 
                           n13687, ZN => n1657);
   U10648 : OAI22_X1 port map( A1 => n14869, A2 => n15146, B1 => n12014, B2 => 
                           n13688, ZN => n1658);
   U10649 : OAI22_X1 port map( A1 => n14869, A2 => n15149, B1 => n12014, B2 => 
                           n13689, ZN => n1659);
   U10650 : OAI22_X1 port map( A1 => n14870, A2 => n15152, B1 => n12014, B2 => 
                           n13690, ZN => n1660);
   U10651 : OAI22_X1 port map( A1 => n14870, A2 => n15164, B1 => n12014, B2 => 
                           n13691, ZN => n1661);
   U10652 : OAI22_X1 port map( A1 => n14877, A2 => n15134, B1 => n12013, B2 => 
                           n13884, ZN => n1686);
   U10653 : OAI22_X1 port map( A1 => n14878, A2 => n15137, B1 => n12013, B2 => 
                           n13885, ZN => n1687);
   U10654 : OAI22_X1 port map( A1 => n14878, A2 => n15140, B1 => n12013, B2 => 
                           n13886, ZN => n1688);
   U10655 : OAI22_X1 port map( A1 => n14878, A2 => n15143, B1 => n12013, B2 => 
                           n13887, ZN => n1689);
   U10656 : OAI22_X1 port map( A1 => n14878, A2 => n15146, B1 => n12013, B2 => 
                           n13888, ZN => n1690);
   U10657 : OAI22_X1 port map( A1 => n14878, A2 => n15149, B1 => n12013, B2 => 
                           n13889, ZN => n1691);
   U10658 : OAI22_X1 port map( A1 => n14879, A2 => n15152, B1 => n12013, B2 => 
                           n13890, ZN => n1692);
   U10659 : OAI22_X1 port map( A1 => n14879, A2 => n15164, B1 => n12013, B2 => 
                           n13891, ZN => n1693);
   U10660 : OAI22_X1 port map( A1 => n14886, A2 => n15134, B1 => n12011, B2 => 
                           n13804, ZN => n1718);
   U10661 : OAI22_X1 port map( A1 => n14887, A2 => n15137, B1 => n12011, B2 => 
                           n13805, ZN => n1719);
   U10662 : OAI22_X1 port map( A1 => n14887, A2 => n15140, B1 => n12011, B2 => 
                           n13806, ZN => n1720);
   U10663 : OAI22_X1 port map( A1 => n14887, A2 => n15143, B1 => n12011, B2 => 
                           n13807, ZN => n1721);
   U10664 : OAI22_X1 port map( A1 => n14887, A2 => n15146, B1 => n12011, B2 => 
                           n13808, ZN => n1722);
   U10665 : OAI22_X1 port map( A1 => n14887, A2 => n15149, B1 => n12011, B2 => 
                           n13809, ZN => n1723);
   U10666 : OAI22_X1 port map( A1 => n14888, A2 => n15152, B1 => n12011, B2 => 
                           n13810, ZN => n1724);
   U10667 : OAI22_X1 port map( A1 => n14888, A2 => n15164, B1 => n12011, B2 => 
                           n13811, ZN => n1725);
   U10668 : OAI22_X1 port map( A1 => n14895, A2 => n15134, B1 => n12009, B2 => 
                           n13893, ZN => n1750);
   U10669 : OAI22_X1 port map( A1 => n14896, A2 => n15137, B1 => n12009, B2 => 
                           n13895, ZN => n1751);
   U10670 : OAI22_X1 port map( A1 => n14896, A2 => n15140, B1 => n12009, B2 => 
                           n13897, ZN => n1752);
   U10671 : OAI22_X1 port map( A1 => n14896, A2 => n15143, B1 => n12009, B2 => 
                           n13899, ZN => n1753);
   U10672 : OAI22_X1 port map( A1 => n14896, A2 => n15146, B1 => n12009, B2 => 
                           n13901, ZN => n1754);
   U10673 : OAI22_X1 port map( A1 => n14896, A2 => n15149, B1 => n12009, B2 => 
                           n13903, ZN => n1755);
   U10674 : OAI22_X1 port map( A1 => n14897, A2 => n15152, B1 => n12009, B2 => 
                           n13905, ZN => n1756);
   U10675 : OAI22_X1 port map( A1 => n14897, A2 => n15164, B1 => n12009, B2 => 
                           n13907, ZN => n1757);
   U10676 : OAI22_X1 port map( A1 => n14904, A2 => n15134, B1 => n12008, B2 => 
                           n13644, ZN => n1782);
   U10677 : OAI22_X1 port map( A1 => n14905, A2 => n15137, B1 => n12008, B2 => 
                           n13645, ZN => n1783);
   U10678 : OAI22_X1 port map( A1 => n14905, A2 => n15140, B1 => n12008, B2 => 
                           n13646, ZN => n1784);
   U10679 : OAI22_X1 port map( A1 => n14905, A2 => n15143, B1 => n12008, B2 => 
                           n13647, ZN => n1785);
   U10680 : OAI22_X1 port map( A1 => n14905, A2 => n15146, B1 => n12008, B2 => 
                           n13648, ZN => n1786);
   U10681 : OAI22_X1 port map( A1 => n14905, A2 => n15149, B1 => n12008, B2 => 
                           n13649, ZN => n1787);
   U10682 : OAI22_X1 port map( A1 => n14906, A2 => n15152, B1 => n12008, B2 => 
                           n13650, ZN => n1788);
   U10683 : OAI22_X1 port map( A1 => n14906, A2 => n15164, B1 => n12008, B2 => 
                           n13651, ZN => n1789);
   U10684 : OAI22_X1 port map( A1 => n14913, A2 => n15134, B1 => n12007, B2 => 
                           n13704, ZN => n1814);
   U10685 : OAI22_X1 port map( A1 => n14914, A2 => n15137, B1 => n12007, B2 => 
                           n13705, ZN => n1815);
   U10686 : OAI22_X1 port map( A1 => n14914, A2 => n15140, B1 => n12007, B2 => 
                           n13706, ZN => n1816);
   U10687 : OAI22_X1 port map( A1 => n14914, A2 => n15143, B1 => n12007, B2 => 
                           n13707, ZN => n1817);
   U10688 : OAI22_X1 port map( A1 => n14914, A2 => n15146, B1 => n12007, B2 => 
                           n13708, ZN => n1818);
   U10689 : OAI22_X1 port map( A1 => n14914, A2 => n15149, B1 => n12007, B2 => 
                           n13709, ZN => n1819);
   U10690 : OAI22_X1 port map( A1 => n14915, A2 => n15152, B1 => n12007, B2 => 
                           n13710, ZN => n1820);
   U10691 : OAI22_X1 port map( A1 => n14915, A2 => n15164, B1 => n12007, B2 => 
                           n13711, ZN => n1821);
   U10692 : OAI22_X1 port map( A1 => n14922, A2 => n15134, B1 => n12005, B2 => 
                           n13872, ZN => n1846);
   U10693 : OAI22_X1 port map( A1 => n14923, A2 => n15137, B1 => n12005, B2 => 
                           n13873, ZN => n1847);
   U10694 : OAI22_X1 port map( A1 => n14923, A2 => n15140, B1 => n12005, B2 => 
                           n13874, ZN => n1848);
   U10695 : OAI22_X1 port map( A1 => n14923, A2 => n15143, B1 => n12005, B2 => 
                           n13875, ZN => n1849);
   U10696 : OAI22_X1 port map( A1 => n14923, A2 => n15146, B1 => n12005, B2 => 
                           n13876, ZN => n1850);
   U10697 : OAI22_X1 port map( A1 => n14923, A2 => n15149, B1 => n12005, B2 => 
                           n13877, ZN => n1851);
   U10698 : OAI22_X1 port map( A1 => n14924, A2 => n15152, B1 => n12005, B2 => 
                           n13878, ZN => n1852);
   U10699 : OAI22_X1 port map( A1 => n14924, A2 => n15164, B1 => n12005, B2 => 
                           n13879, ZN => n1853);
   U10700 : OAI22_X1 port map( A1 => n14976, A2 => n15133, B1 => n11998, B2 => 
                           n13652, ZN => n2038);
   U10701 : OAI22_X1 port map( A1 => n14977, A2 => n15136, B1 => n11998, B2 => 
                           n13653, ZN => n2039);
   U10702 : OAI22_X1 port map( A1 => n14977, A2 => n15139, B1 => n11998, B2 => 
                           n13654, ZN => n2040);
   U10703 : OAI22_X1 port map( A1 => n14977, A2 => n15142, B1 => n11998, B2 => 
                           n13655, ZN => n2041);
   U10704 : OAI22_X1 port map( A1 => n14977, A2 => n15145, B1 => n11998, B2 => 
                           n13656, ZN => n2042);
   U10705 : OAI22_X1 port map( A1 => n14977, A2 => n15148, B1 => n11998, B2 => 
                           n13657, ZN => n2043);
   U10706 : OAI22_X1 port map( A1 => n14978, A2 => n15151, B1 => n11998, B2 => 
                           n13658, ZN => n2044);
   U10707 : OAI22_X1 port map( A1 => n14978, A2 => n15163, B1 => n11998, B2 => 
                           n13659, ZN => n2045);
   U10708 : OAI22_X1 port map( A1 => n14985, A2 => n15133, B1 => n11997, B2 => 
                           n13856, ZN => n2070);
   U10709 : OAI22_X1 port map( A1 => n14986, A2 => n15136, B1 => n11997, B2 => 
                           n13857, ZN => n2071);
   U10710 : OAI22_X1 port map( A1 => n14986, A2 => n15139, B1 => n11997, B2 => 
                           n13858, ZN => n2072);
   U10711 : OAI22_X1 port map( A1 => n14986, A2 => n15142, B1 => n11997, B2 => 
                           n13859, ZN => n2073);
   U10712 : OAI22_X1 port map( A1 => n14986, A2 => n15145, B1 => n11997, B2 => 
                           n13860, ZN => n2074);
   U10713 : OAI22_X1 port map( A1 => n14986, A2 => n15148, B1 => n11997, B2 => 
                           n13861, ZN => n2075);
   U10714 : OAI22_X1 port map( A1 => n14987, A2 => n15151, B1 => n11997, B2 => 
                           n13862, ZN => n2076);
   U10715 : OAI22_X1 port map( A1 => n14987, A2 => n15163, B1 => n11997, B2 => 
                           n13863, ZN => n2077);
   U10716 : OAI22_X1 port map( A1 => n14994, A2 => n15133, B1 => n11995, B2 => 
                           n13752, ZN => n2102);
   U10717 : OAI22_X1 port map( A1 => n14995, A2 => n15136, B1 => n11995, B2 => 
                           n13753, ZN => n2103);
   U10718 : OAI22_X1 port map( A1 => n14995, A2 => n15139, B1 => n11995, B2 => 
                           n13754, ZN => n2104);
   U10719 : OAI22_X1 port map( A1 => n14995, A2 => n15142, B1 => n11995, B2 => 
                           n13755, ZN => n2105);
   U10720 : OAI22_X1 port map( A1 => n14995, A2 => n15145, B1 => n11995, B2 => 
                           n13756, ZN => n2106);
   U10721 : OAI22_X1 port map( A1 => n14995, A2 => n15148, B1 => n11995, B2 => 
                           n13757, ZN => n2107);
   U10722 : OAI22_X1 port map( A1 => n14996, A2 => n15151, B1 => n11995, B2 => 
                           n13758, ZN => n2108);
   U10723 : OAI22_X1 port map( A1 => n14996, A2 => n15163, B1 => n11995, B2 => 
                           n13759, ZN => n2109);
   U10724 : OAI22_X1 port map( A1 => n15048, A2 => n15133, B1 => n11985, B2 => 
                           n13824, ZN => n2294);
   U10725 : OAI22_X1 port map( A1 => n15049, A2 => n15136, B1 => n11985, B2 => 
                           n13825, ZN => n2295);
   U10726 : OAI22_X1 port map( A1 => n15049, A2 => n15139, B1 => n11985, B2 => 
                           n13826, ZN => n2296);
   U10727 : OAI22_X1 port map( A1 => n15049, A2 => n15142, B1 => n11985, B2 => 
                           n13827, ZN => n2297);
   U10728 : OAI22_X1 port map( A1 => n15049, A2 => n15145, B1 => n11985, B2 => 
                           n13828, ZN => n2298);
   U10729 : OAI22_X1 port map( A1 => n15049, A2 => n15148, B1 => n11985, B2 => 
                           n13829, ZN => n2299);
   U10730 : OAI22_X1 port map( A1 => n15050, A2 => n15151, B1 => n11985, B2 => 
                           n13830, ZN => n2300);
   U10731 : OAI22_X1 port map( A1 => n15050, A2 => n15163, B1 => n11985, B2 => 
                           n13831, ZN => n2301);
   U10732 : OAI22_X1 port map( A1 => n15057, A2 => n15133, B1 => n11983, B2 => 
                           n13864, ZN => n2326);
   U10733 : OAI22_X1 port map( A1 => n15058, A2 => n15136, B1 => n11983, B2 => 
                           n13865, ZN => n2327);
   U10734 : OAI22_X1 port map( A1 => n15058, A2 => n15139, B1 => n11983, B2 => 
                           n13866, ZN => n2328);
   U10735 : OAI22_X1 port map( A1 => n15058, A2 => n15142, B1 => n11983, B2 => 
                           n13867, ZN => n2329);
   U10736 : OAI22_X1 port map( A1 => n15058, A2 => n15145, B1 => n11983, B2 => 
                           n13868, ZN => n2330);
   U10737 : OAI22_X1 port map( A1 => n15058, A2 => n15148, B1 => n11983, B2 => 
                           n13869, ZN => n2331);
   U10738 : OAI22_X1 port map( A1 => n15059, A2 => n15151, B1 => n11983, B2 => 
                           n13870, ZN => n2332);
   U10739 : OAI22_X1 port map( A1 => n15059, A2 => n15163, B1 => n11983, B2 => 
                           n13871, ZN => n2333);
   U10740 : OAI22_X1 port map( A1 => n15159, A2 => n15133, B1 => n11949, B2 => 
                           n13760, ZN => n2358);
   U10741 : OAI22_X1 port map( A1 => n15160, A2 => n15136, B1 => n11949, B2 => 
                           n13761, ZN => n2359);
   U10742 : OAI22_X1 port map( A1 => n15160, A2 => n15139, B1 => n11949, B2 => 
                           n13762, ZN => n2360);
   U10743 : OAI22_X1 port map( A1 => n15160, A2 => n15142, B1 => n11949, B2 => 
                           n13763, ZN => n2361);
   U10744 : OAI22_X1 port map( A1 => n15160, A2 => n15145, B1 => n11949, B2 => 
                           n13764, ZN => n2362);
   U10745 : OAI22_X1 port map( A1 => n15160, A2 => n15148, B1 => n11949, B2 => 
                           n13765, ZN => n2363);
   U10746 : OAI22_X1 port map( A1 => n15161, A2 => n15151, B1 => n11949, B2 => 
                           n13766, ZN => n2364);
   U10747 : OAI22_X1 port map( A1 => n15161, A2 => n15163, B1 => n11949, B2 => 
                           n13767, ZN => n2365);
   U10748 : AOI22_X1 port map( A1 => n14626, A2 => n13916, B1 => n14625, B2 => 
                           n14322, ZN => n13184);
   U10749 : AOI22_X1 port map( A1 => n14626, A2 => n13917, B1 => n14625, B2 => 
                           n14323, ZN => n13164);
   U10750 : AOI22_X1 port map( A1 => n14626, A2 => n13918, B1 => n14625, B2 => 
                           n14324, ZN => n13147);
   U10751 : AOI22_X1 port map( A1 => n14626, A2 => n13919, B1 => n14625, B2 => 
                           n14325, ZN => n13130);
   U10752 : AOI22_X1 port map( A1 => n14626, A2 => n13920, B1 => n14625, B2 => 
                           n14326, ZN => n13113);
   U10753 : AOI22_X1 port map( A1 => n14626, A2 => n13921, B1 => n14625, B2 => 
                           n14327, ZN => n13096);
   U10754 : AOI22_X1 port map( A1 => n14626, A2 => n13922, B1 => n14625, B2 => 
                           n14328, ZN => n13079);
   U10755 : AOI22_X1 port map( A1 => n14626, A2 => n13923, B1 => n14625, B2 => 
                           n14329, ZN => n13062);
   U10756 : AOI22_X1 port map( A1 => n14626, A2 => n13924, B1 => n14624, B2 => 
                           n14330, ZN => n13045);
   U10757 : AOI22_X1 port map( A1 => n14626, A2 => n13925, B1 => n14624, B2 => 
                           n14331, ZN => n13028);
   U10758 : AOI22_X1 port map( A1 => n14626, A2 => n13926, B1 => n14624, B2 => 
                           n14332, ZN => n13011);
   U10759 : AOI22_X1 port map( A1 => n14626, A2 => n13927, B1 => n14624, B2 => 
                           n14333, ZN => n12994);
   U10760 : AOI22_X1 port map( A1 => n14627, A2 => n13928, B1 => n14624, B2 => 
                           n14334, ZN => n12977);
   U10761 : AOI22_X1 port map( A1 => n14627, A2 => n13929, B1 => n14624, B2 => 
                           n14335, ZN => n12960);
   U10762 : AOI22_X1 port map( A1 => n14627, A2 => n13930, B1 => n14624, B2 => 
                           n14336, ZN => n12943);
   U10763 : AOI22_X1 port map( A1 => n14627, A2 => n13931, B1 => n14624, B2 => 
                           n14337, ZN => n12926);
   U10764 : AOI22_X1 port map( A1 => n14627, A2 => n13932, B1 => n14624, B2 => 
                           n14338, ZN => n12909);
   U10765 : AOI22_X1 port map( A1 => n14627, A2 => n13933, B1 => n14624, B2 => 
                           n14339, ZN => n12892);
   U10766 : AOI22_X1 port map( A1 => n14627, A2 => n13934, B1 => n14624, B2 => 
                           n14340, ZN => n12875);
   U10767 : AOI22_X1 port map( A1 => n14627, A2 => n13935, B1 => n14624, B2 => 
                           n14341, ZN => n12858);
   U10768 : AOI22_X1 port map( A1 => n14627, A2 => n13936, B1 => n14623, B2 => 
                           n14342, ZN => n12841);
   U10769 : AOI22_X1 port map( A1 => n14627, A2 => n13937, B1 => n14623, B2 => 
                           n14343, ZN => n12824);
   U10770 : AOI22_X1 port map( A1 => n14627, A2 => n13938, B1 => n14623, B2 => 
                           n14344, ZN => n12807);
   U10771 : AOI22_X1 port map( A1 => n14627, A2 => n13939, B1 => n14623, B2 => 
                           n14345, ZN => n12790);
   U10772 : AOI22_X1 port map( A1 => n14628, A2 => n13940, B1 => n14623, B2 => 
                           n14346, ZN => n12773);
   U10773 : AOI22_X1 port map( A1 => n14628, A2 => n13941, B1 => n14623, B2 => 
                           n14347, ZN => n12756);
   U10774 : AOI22_X1 port map( A1 => n14628, A2 => n13942, B1 => n14623, B2 => 
                           n14348, ZN => n12739);
   U10775 : AOI22_X1 port map( A1 => n14628, A2 => n13943, B1 => n14623, B2 => 
                           n14349, ZN => n12722);
   U10776 : AOI22_X1 port map( A1 => n14628, A2 => n13944, B1 => n14623, B2 => 
                           n14350, ZN => n12705);
   U10777 : AOI22_X1 port map( A1 => n14628, A2 => n13945, B1 => n14623, B2 => 
                           n14351, ZN => n12688);
   U10778 : AOI22_X1 port map( A1 => n14628, A2 => n13946, B1 => n14623, B2 => 
                           n14352, ZN => n12671);
   U10779 : AOI22_X1 port map( A1 => n14628, A2 => n13947, B1 => n14623, B2 => 
                           n14353, ZN => n12639);
   U10780 : AOI22_X1 port map( A1 => n14724, A2 => n13916, B1 => n14723, B2 => 
                           n14322, ZN => n12603);
   U10781 : AOI22_X1 port map( A1 => n14724, A2 => n13917, B1 => n14723, B2 => 
                           n14323, ZN => n12583);
   U10782 : AOI22_X1 port map( A1 => n14724, A2 => n13918, B1 => n14723, B2 => 
                           n14324, ZN => n12566);
   U10783 : AOI22_X1 port map( A1 => n14724, A2 => n13919, B1 => n14723, B2 => 
                           n14325, ZN => n12549);
   U10784 : AOI22_X1 port map( A1 => n14724, A2 => n13920, B1 => n14723, B2 => 
                           n14326, ZN => n12532);
   U10785 : AOI22_X1 port map( A1 => n14724, A2 => n13921, B1 => n14723, B2 => 
                           n14327, ZN => n12515);
   U10786 : AOI22_X1 port map( A1 => n14724, A2 => n13922, B1 => n14723, B2 => 
                           n14328, ZN => n12498);
   U10787 : AOI22_X1 port map( A1 => n14724, A2 => n13923, B1 => n14723, B2 => 
                           n14329, ZN => n12481);
   U10788 : AOI22_X1 port map( A1 => n14724, A2 => n13924, B1 => n14722, B2 => 
                           n14330, ZN => n12464);
   U10789 : AOI22_X1 port map( A1 => n14724, A2 => n13925, B1 => n14722, B2 => 
                           n14331, ZN => n12447);
   U10790 : AOI22_X1 port map( A1 => n14724, A2 => n13926, B1 => n14722, B2 => 
                           n14332, ZN => n12430);
   U10791 : AOI22_X1 port map( A1 => n14724, A2 => n13927, B1 => n14722, B2 => 
                           n14333, ZN => n12413);
   U10792 : AOI22_X1 port map( A1 => n14725, A2 => n13928, B1 => n14722, B2 => 
                           n14334, ZN => n12396);
   U10793 : AOI22_X1 port map( A1 => n14725, A2 => n13929, B1 => n14722, B2 => 
                           n14335, ZN => n12379);
   U10794 : AOI22_X1 port map( A1 => n14725, A2 => n13930, B1 => n14722, B2 => 
                           n14336, ZN => n12362);
   U10795 : AOI22_X1 port map( A1 => n14725, A2 => n13931, B1 => n14722, B2 => 
                           n14337, ZN => n12345);
   U10796 : AOI22_X1 port map( A1 => n14725, A2 => n13932, B1 => n14722, B2 => 
                           n14338, ZN => n12328);
   U10797 : AOI22_X1 port map( A1 => n14725, A2 => n13933, B1 => n14722, B2 => 
                           n14339, ZN => n12311);
   U10798 : AOI22_X1 port map( A1 => n14725, A2 => n13934, B1 => n14722, B2 => 
                           n14340, ZN => n12294);
   U10799 : AOI22_X1 port map( A1 => n14725, A2 => n13935, B1 => n14722, B2 => 
                           n14341, ZN => n12277);
   U10800 : AOI22_X1 port map( A1 => n14725, A2 => n13936, B1 => n14721, B2 => 
                           n14342, ZN => n12260);
   U10801 : AOI22_X1 port map( A1 => n14725, A2 => n13937, B1 => n14721, B2 => 
                           n14343, ZN => n12243);
   U10802 : AOI22_X1 port map( A1 => n14725, A2 => n13938, B1 => n14721, B2 => 
                           n14344, ZN => n12226);
   U10803 : AOI22_X1 port map( A1 => n14725, A2 => n13939, B1 => n14721, B2 => 
                           n14345, ZN => n12209);
   U10804 : AOI22_X1 port map( A1 => n14726, A2 => n13940, B1 => n14721, B2 => 
                           n14346, ZN => n12192);
   U10805 : AOI22_X1 port map( A1 => n14726, A2 => n13941, B1 => n14721, B2 => 
                           n14347, ZN => n12175);
   U10806 : AOI22_X1 port map( A1 => n14726, A2 => n13942, B1 => n14721, B2 => 
                           n14348, ZN => n12158);
   U10807 : AOI22_X1 port map( A1 => n14726, A2 => n13943, B1 => n14721, B2 => 
                           n14349, ZN => n12141);
   U10808 : AOI22_X1 port map( A1 => n14726, A2 => n13944, B1 => n14721, B2 => 
                           n14350, ZN => n12124);
   U10809 : AOI22_X1 port map( A1 => n14726, A2 => n13945, B1 => n14721, B2 => 
                           n14351, ZN => n12107);
   U10810 : AOI22_X1 port map( A1 => n14726, A2 => n13946, B1 => n14721, B2 => 
                           n14352, ZN => n12090);
   U10811 : AOI22_X1 port map( A1 => n14726, A2 => n13947, B1 => n14721, B2 => 
                           n14353, ZN => n12058);
   U10812 : OAI22_X1 port map( A1 => n14855, A2 => n15062, B1 => n14854, B2 => 
                           n13908, ZN => n1598);
   U10813 : OAI22_X1 port map( A1 => n14855, A2 => n15065, B1 => n14854, B2 => 
                           n13909, ZN => n1599);
   U10814 : OAI22_X1 port map( A1 => n14855, A2 => n15068, B1 => n14854, B2 => 
                           n13910, ZN => n1600);
   U10815 : OAI22_X1 port map( A1 => n14855, A2 => n15071, B1 => n14854, B2 => 
                           n13911, ZN => n1601);
   U10816 : OAI22_X1 port map( A1 => n14855, A2 => n15074, B1 => n14854, B2 => 
                           n13912, ZN => n1602);
   U10817 : OAI22_X1 port map( A1 => n14856, A2 => n15077, B1 => n14854, B2 => 
                           n13913, ZN => n1603);
   U10818 : OAI22_X1 port map( A1 => n14856, A2 => n15080, B1 => n14854, B2 => 
                           n13914, ZN => n1604);
   U10819 : OAI22_X1 port map( A1 => n14856, A2 => n15083, B1 => n14854, B2 => 
                           n13915, ZN => n1605);
   U10820 : OAI22_X1 port map( A1 => n14856, A2 => n15086, B1 => n14854, B2 => 
                           n13880, ZN => n1606);
   U10821 : OAI22_X1 port map( A1 => n14856, A2 => n15089, B1 => n14854, B2 => 
                           n13881, ZN => n1607);
   U10822 : OAI22_X1 port map( A1 => n14857, A2 => n15092, B1 => n14854, B2 => 
                           n13882, ZN => n1608);
   U10823 : OAI22_X1 port map( A1 => n14857, A2 => n15095, B1 => n14854, B2 => 
                           n13883, ZN => n1609);
   U10824 : OAI22_X1 port map( A1 => n14857, A2 => n15098, B1 => n12015, B2 => 
                           n14170, ZN => n1610);
   U10825 : OAI22_X1 port map( A1 => n14857, A2 => n15101, B1 => n12015, B2 => 
                           n14172, ZN => n1611);
   U10826 : OAI22_X1 port map( A1 => n14857, A2 => n15104, B1 => n12015, B2 => 
                           n14174, ZN => n1612);
   U10827 : OAI22_X1 port map( A1 => n14858, A2 => n15107, B1 => n14854, B2 => 
                           n14176, ZN => n1613);
   U10828 : OAI22_X1 port map( A1 => n14858, A2 => n15110, B1 => n14854, B2 => 
                           n14178, ZN => n1614);
   U10829 : OAI22_X1 port map( A1 => n14858, A2 => n15113, B1 => n14854, B2 => 
                           n14180, ZN => n1615);
   U10830 : OAI22_X1 port map( A1 => n14858, A2 => n15116, B1 => n14854, B2 => 
                           n14182, ZN => n1616);
   U10831 : OAI22_X1 port map( A1 => n14858, A2 => n15119, B1 => n14854, B2 => 
                           n14184, ZN => n1617);
   U10832 : OAI22_X1 port map( A1 => n14859, A2 => n15122, B1 => n14854, B2 => 
                           n14186, ZN => n1618);
   U10833 : OAI22_X1 port map( A1 => n14859, A2 => n15125, B1 => n14854, B2 => 
                           n14188, ZN => n1619);
   U10834 : OAI22_X1 port map( A1 => n14859, A2 => n15128, B1 => n14854, B2 => 
                           n14190, ZN => n1620);
   U10835 : OAI22_X1 port map( A1 => n14859, A2 => n15131, B1 => n14854, B2 => 
                           n14192, ZN => n1621);
   U10836 : OAI22_X1 port map( A1 => n14864, A2 => n15062, B1 => n14863, B2 => 
                           n13792, ZN => n1630);
   U10837 : OAI22_X1 port map( A1 => n14864, A2 => n15065, B1 => n14863, B2 => 
                           n13793, ZN => n1631);
   U10838 : OAI22_X1 port map( A1 => n14864, A2 => n15068, B1 => n14863, B2 => 
                           n13794, ZN => n1632);
   U10839 : OAI22_X1 port map( A1 => n14864, A2 => n15071, B1 => n14863, B2 => 
                           n13795, ZN => n1633);
   U10840 : OAI22_X1 port map( A1 => n14864, A2 => n15074, B1 => n14863, B2 => 
                           n13796, ZN => n1634);
   U10841 : OAI22_X1 port map( A1 => n14865, A2 => n15077, B1 => n14863, B2 => 
                           n13797, ZN => n1635);
   U10842 : OAI22_X1 port map( A1 => n14865, A2 => n15080, B1 => n14863, B2 => 
                           n13798, ZN => n1636);
   U10843 : OAI22_X1 port map( A1 => n14865, A2 => n15083, B1 => n14863, B2 => 
                           n13799, ZN => n1637);
   U10844 : OAI22_X1 port map( A1 => n14865, A2 => n15086, B1 => n14863, B2 => 
                           n13800, ZN => n1638);
   U10845 : OAI22_X1 port map( A1 => n14865, A2 => n15089, B1 => n14863, B2 => 
                           n13801, ZN => n1639);
   U10846 : OAI22_X1 port map( A1 => n14866, A2 => n15092, B1 => n14863, B2 => 
                           n13802, ZN => n1640);
   U10847 : OAI22_X1 port map( A1 => n14866, A2 => n15095, B1 => n14863, B2 => 
                           n13803, ZN => n1641);
   U10848 : OAI22_X1 port map( A1 => n14866, A2 => n15098, B1 => n12014, B2 => 
                           n13692, ZN => n1642);
   U10849 : OAI22_X1 port map( A1 => n14866, A2 => n15101, B1 => n12014, B2 => 
                           n13693, ZN => n1643);
   U10850 : OAI22_X1 port map( A1 => n14866, A2 => n15104, B1 => n12014, B2 => 
                           n13694, ZN => n1644);
   U10851 : OAI22_X1 port map( A1 => n14867, A2 => n15107, B1 => n14863, B2 => 
                           n13695, ZN => n1645);
   U10852 : OAI22_X1 port map( A1 => n14867, A2 => n15110, B1 => n14863, B2 => 
                           n13696, ZN => n1646);
   U10853 : OAI22_X1 port map( A1 => n14867, A2 => n15113, B1 => n14863, B2 => 
                           n13697, ZN => n1647);
   U10854 : OAI22_X1 port map( A1 => n14867, A2 => n15116, B1 => n14863, B2 => 
                           n13698, ZN => n1648);
   U10855 : OAI22_X1 port map( A1 => n14867, A2 => n15119, B1 => n14863, B2 => 
                           n13699, ZN => n1649);
   U10856 : OAI22_X1 port map( A1 => n14868, A2 => n15122, B1 => n14863, B2 => 
                           n13700, ZN => n1650);
   U10857 : OAI22_X1 port map( A1 => n14868, A2 => n15125, B1 => n14863, B2 => 
                           n13701, ZN => n1651);
   U10858 : OAI22_X1 port map( A1 => n14868, A2 => n15128, B1 => n14863, B2 => 
                           n13702, ZN => n1652);
   U10859 : OAI22_X1 port map( A1 => n14868, A2 => n15131, B1 => n14863, B2 => 
                           n13703, ZN => n1653);
   U10860 : OAI22_X1 port map( A1 => n14873, A2 => n15062, B1 => n14872, B2 => 
                           n14194, ZN => n1662);
   U10861 : OAI22_X1 port map( A1 => n14873, A2 => n15065, B1 => n14872, B2 => 
                           n14195, ZN => n1663);
   U10862 : OAI22_X1 port map( A1 => n14873, A2 => n15068, B1 => n14872, B2 => 
                           n14196, ZN => n1664);
   U10863 : OAI22_X1 port map( A1 => n14873, A2 => n15071, B1 => n14872, B2 => 
                           n14197, ZN => n1665);
   U10864 : OAI22_X1 port map( A1 => n14873, A2 => n15074, B1 => n14872, B2 => 
                           n14198, ZN => n1666);
   U10865 : OAI22_X1 port map( A1 => n14874, A2 => n15077, B1 => n14872, B2 => 
                           n14199, ZN => n1667);
   U10866 : OAI22_X1 port map( A1 => n14874, A2 => n15080, B1 => n14872, B2 => 
                           n14200, ZN => n1668);
   U10867 : OAI22_X1 port map( A1 => n14874, A2 => n15083, B1 => n14872, B2 => 
                           n14201, ZN => n1669);
   U10868 : OAI22_X1 port map( A1 => n14874, A2 => n15086, B1 => n14872, B2 => 
                           n14202, ZN => n1670);
   U10869 : OAI22_X1 port map( A1 => n14874, A2 => n15089, B1 => n14872, B2 => 
                           n14203, ZN => n1671);
   U10870 : OAI22_X1 port map( A1 => n14875, A2 => n15092, B1 => n14872, B2 => 
                           n14204, ZN => n1672);
   U10871 : OAI22_X1 port map( A1 => n14875, A2 => n15095, B1 => n14872, B2 => 
                           n14205, ZN => n1673);
   U10872 : OAI22_X1 port map( A1 => n14875, A2 => n15098, B1 => n12013, B2 => 
                           n14206, ZN => n1674);
   U10873 : OAI22_X1 port map( A1 => n14875, A2 => n15101, B1 => n12013, B2 => 
                           n14207, ZN => n1675);
   U10874 : OAI22_X1 port map( A1 => n14875, A2 => n15104, B1 => n12013, B2 => 
                           n14208, ZN => n1676);
   U10875 : OAI22_X1 port map( A1 => n14876, A2 => n15107, B1 => n14872, B2 => 
                           n14209, ZN => n1677);
   U10876 : OAI22_X1 port map( A1 => n14876, A2 => n15110, B1 => n14872, B2 => 
                           n14210, ZN => n1678);
   U10877 : OAI22_X1 port map( A1 => n14876, A2 => n15113, B1 => n14872, B2 => 
                           n14211, ZN => n1679);
   U10878 : OAI22_X1 port map( A1 => n14876, A2 => n15116, B1 => n14872, B2 => 
                           n14212, ZN => n1680);
   U10879 : OAI22_X1 port map( A1 => n14876, A2 => n15119, B1 => n14872, B2 => 
                           n14213, ZN => n1681);
   U10880 : OAI22_X1 port map( A1 => n14877, A2 => n15122, B1 => n14872, B2 => 
                           n14214, ZN => n1682);
   U10881 : OAI22_X1 port map( A1 => n14877, A2 => n15125, B1 => n14872, B2 => 
                           n14215, ZN => n1683);
   U10882 : OAI22_X1 port map( A1 => n14877, A2 => n15128, B1 => n14872, B2 => 
                           n14216, ZN => n1684);
   U10883 : OAI22_X1 port map( A1 => n14877, A2 => n15131, B1 => n14872, B2 => 
                           n14217, ZN => n1685);
   U10884 : OAI22_X1 port map( A1 => n14882, A2 => n15062, B1 => n14881, B2 => 
                           n14046, ZN => n1694);
   U10885 : OAI22_X1 port map( A1 => n14882, A2 => n15065, B1 => n14881, B2 => 
                           n14047, ZN => n1695);
   U10886 : OAI22_X1 port map( A1 => n14882, A2 => n15068, B1 => n14881, B2 => 
                           n14048, ZN => n1696);
   U10887 : OAI22_X1 port map( A1 => n14882, A2 => n15071, B1 => n14881, B2 => 
                           n14049, ZN => n1697);
   U10888 : OAI22_X1 port map( A1 => n14882, A2 => n15074, B1 => n14881, B2 => 
                           n14050, ZN => n1698);
   U10889 : OAI22_X1 port map( A1 => n14883, A2 => n15077, B1 => n14881, B2 => 
                           n14051, ZN => n1699);
   U10890 : OAI22_X1 port map( A1 => n14883, A2 => n15080, B1 => n14881, B2 => 
                           n14052, ZN => n1700);
   U10891 : OAI22_X1 port map( A1 => n14883, A2 => n15083, B1 => n14881, B2 => 
                           n14053, ZN => n1701);
   U10892 : OAI22_X1 port map( A1 => n14883, A2 => n15086, B1 => n14881, B2 => 
                           n14054, ZN => n1702);
   U10893 : OAI22_X1 port map( A1 => n14883, A2 => n15089, B1 => n14881, B2 => 
                           n14055, ZN => n1703);
   U10894 : OAI22_X1 port map( A1 => n14884, A2 => n15092, B1 => n14881, B2 => 
                           n14056, ZN => n1704);
   U10895 : OAI22_X1 port map( A1 => n14884, A2 => n15095, B1 => n14881, B2 => 
                           n14057, ZN => n1705);
   U10896 : OAI22_X1 port map( A1 => n14884, A2 => n15098, B1 => n12011, B2 => 
                           n14058, ZN => n1706);
   U10897 : OAI22_X1 port map( A1 => n14884, A2 => n15101, B1 => n12011, B2 => 
                           n14059, ZN => n1707);
   U10898 : OAI22_X1 port map( A1 => n14884, A2 => n15104, B1 => n12011, B2 => 
                           n14060, ZN => n1708);
   U10899 : OAI22_X1 port map( A1 => n14885, A2 => n15107, B1 => n14881, B2 => 
                           n14061, ZN => n1709);
   U10900 : OAI22_X1 port map( A1 => n14885, A2 => n15110, B1 => n14881, B2 => 
                           n14062, ZN => n1710);
   U10901 : OAI22_X1 port map( A1 => n14885, A2 => n15113, B1 => n14881, B2 => 
                           n14063, ZN => n1711);
   U10902 : OAI22_X1 port map( A1 => n14885, A2 => n15116, B1 => n14881, B2 => 
                           n14064, ZN => n1712);
   U10903 : OAI22_X1 port map( A1 => n14885, A2 => n15119, B1 => n14881, B2 => 
                           n14065, ZN => n1713);
   U10904 : OAI22_X1 port map( A1 => n14886, A2 => n15122, B1 => n14881, B2 => 
                           n14066, ZN => n1714);
   U10905 : OAI22_X1 port map( A1 => n14886, A2 => n15125, B1 => n14881, B2 => 
                           n14067, ZN => n1715);
   U10906 : OAI22_X1 port map( A1 => n14886, A2 => n15128, B1 => n14881, B2 => 
                           n14068, ZN => n1716);
   U10907 : OAI22_X1 port map( A1 => n14886, A2 => n15131, B1 => n14881, B2 => 
                           n14069, ZN => n1717);
   U10908 : OAI22_X1 port map( A1 => n14891, A2 => n15062, B1 => n14890, B2 => 
                           n14218, ZN => n1726);
   U10909 : OAI22_X1 port map( A1 => n14891, A2 => n15065, B1 => n14890, B2 => 
                           n14219, ZN => n1727);
   U10910 : OAI22_X1 port map( A1 => n14891, A2 => n15068, B1 => n14890, B2 => 
                           n14220, ZN => n1728);
   U10911 : OAI22_X1 port map( A1 => n14891, A2 => n15071, B1 => n14890, B2 => 
                           n14221, ZN => n1729);
   U10912 : OAI22_X1 port map( A1 => n14891, A2 => n15074, B1 => n14890, B2 => 
                           n14222, ZN => n1730);
   U10913 : OAI22_X1 port map( A1 => n14892, A2 => n15077, B1 => n14890, B2 => 
                           n14223, ZN => n1731);
   U10914 : OAI22_X1 port map( A1 => n14892, A2 => n15080, B1 => n14890, B2 => 
                           n14224, ZN => n1732);
   U10915 : OAI22_X1 port map( A1 => n14892, A2 => n15083, B1 => n14890, B2 => 
                           n14225, ZN => n1733);
   U10916 : OAI22_X1 port map( A1 => n14892, A2 => n15086, B1 => n14890, B2 => 
                           n14166, ZN => n1734);
   U10917 : OAI22_X1 port map( A1 => n14892, A2 => n15089, B1 => n14890, B2 => 
                           n14167, ZN => n1735);
   U10918 : OAI22_X1 port map( A1 => n14893, A2 => n15092, B1 => n14890, B2 => 
                           n14168, ZN => n1736);
   U10919 : OAI22_X1 port map( A1 => n14893, A2 => n15095, B1 => n14890, B2 => 
                           n14169, ZN => n1737);
   U10920 : OAI22_X1 port map( A1 => n14893, A2 => n15098, B1 => n12009, B2 => 
                           n14171, ZN => n1738);
   U10921 : OAI22_X1 port map( A1 => n14893, A2 => n15101, B1 => n12009, B2 => 
                           n14173, ZN => n1739);
   U10922 : OAI22_X1 port map( A1 => n14893, A2 => n15104, B1 => n12009, B2 => 
                           n14175, ZN => n1740);
   U10923 : OAI22_X1 port map( A1 => n14894, A2 => n15107, B1 => n14890, B2 => 
                           n14177, ZN => n1741);
   U10924 : OAI22_X1 port map( A1 => n14894, A2 => n15110, B1 => n14890, B2 => 
                           n14179, ZN => n1742);
   U10925 : OAI22_X1 port map( A1 => n14894, A2 => n15113, B1 => n14890, B2 => 
                           n14181, ZN => n1743);
   U10926 : OAI22_X1 port map( A1 => n14894, A2 => n15116, B1 => n14890, B2 => 
                           n14183, ZN => n1744);
   U10927 : OAI22_X1 port map( A1 => n14894, A2 => n15119, B1 => n14890, B2 => 
                           n14185, ZN => n1745);
   U10928 : OAI22_X1 port map( A1 => n14895, A2 => n15122, B1 => n14890, B2 => 
                           n14187, ZN => n1746);
   U10929 : OAI22_X1 port map( A1 => n14895, A2 => n15125, B1 => n14890, B2 => 
                           n14189, ZN => n1747);
   U10930 : OAI22_X1 port map( A1 => n14895, A2 => n15128, B1 => n14890, B2 => 
                           n14191, ZN => n1748);
   U10931 : OAI22_X1 port map( A1 => n14895, A2 => n15131, B1 => n14890, B2 => 
                           n14193, ZN => n1749);
   U10932 : OAI22_X1 port map( A1 => n14900, A2 => n15062, B1 => n14899, B2 => 
                           n13728, ZN => n1758);
   U10933 : OAI22_X1 port map( A1 => n14900, A2 => n15065, B1 => n14899, B2 => 
                           n13729, ZN => n1759);
   U10934 : OAI22_X1 port map( A1 => n14900, A2 => n15068, B1 => n14899, B2 => 
                           n13730, ZN => n1760);
   U10935 : OAI22_X1 port map( A1 => n14900, A2 => n15071, B1 => n14899, B2 => 
                           n13731, ZN => n1761);
   U10936 : OAI22_X1 port map( A1 => n14900, A2 => n15074, B1 => n14899, B2 => 
                           n13732, ZN => n1762);
   U10937 : OAI22_X1 port map( A1 => n14901, A2 => n15077, B1 => n14899, B2 => 
                           n13733, ZN => n1763);
   U10938 : OAI22_X1 port map( A1 => n14901, A2 => n15080, B1 => n14899, B2 => 
                           n13734, ZN => n1764);
   U10939 : OAI22_X1 port map( A1 => n14901, A2 => n15083, B1 => n14899, B2 => 
                           n13735, ZN => n1765);
   U10940 : OAI22_X1 port map( A1 => n14901, A2 => n15086, B1 => n14899, B2 => 
                           n13736, ZN => n1766);
   U10941 : OAI22_X1 port map( A1 => n14901, A2 => n15089, B1 => n14899, B2 => 
                           n13737, ZN => n1767);
   U10942 : OAI22_X1 port map( A1 => n14902, A2 => n15092, B1 => n14899, B2 => 
                           n13738, ZN => n1768);
   U10943 : OAI22_X1 port map( A1 => n14902, A2 => n15095, B1 => n14899, B2 => 
                           n13739, ZN => n1769);
   U10944 : OAI22_X1 port map( A1 => n14902, A2 => n15098, B1 => n12008, B2 => 
                           n13660, ZN => n1770);
   U10945 : OAI22_X1 port map( A1 => n14902, A2 => n15101, B1 => n12008, B2 => 
                           n13661, ZN => n1771);
   U10946 : OAI22_X1 port map( A1 => n14902, A2 => n15104, B1 => n12008, B2 => 
                           n13662, ZN => n1772);
   U10947 : OAI22_X1 port map( A1 => n14903, A2 => n15107, B1 => n14899, B2 => 
                           n13663, ZN => n1773);
   U10948 : OAI22_X1 port map( A1 => n14903, A2 => n15110, B1 => n14899, B2 => 
                           n13664, ZN => n1774);
   U10949 : OAI22_X1 port map( A1 => n14903, A2 => n15113, B1 => n14899, B2 => 
                           n13665, ZN => n1775);
   U10950 : OAI22_X1 port map( A1 => n14903, A2 => n15116, B1 => n14899, B2 => 
                           n13666, ZN => n1776);
   U10951 : OAI22_X1 port map( A1 => n14903, A2 => n15119, B1 => n14899, B2 => 
                           n13667, ZN => n1777);
   U10952 : OAI22_X1 port map( A1 => n14904, A2 => n15122, B1 => n14899, B2 => 
                           n13668, ZN => n1778);
   U10953 : OAI22_X1 port map( A1 => n14904, A2 => n15125, B1 => n14899, B2 => 
                           n13669, ZN => n1779);
   U10954 : OAI22_X1 port map( A1 => n14904, A2 => n15128, B1 => n14899, B2 => 
                           n13670, ZN => n1780);
   U10955 : OAI22_X1 port map( A1 => n14904, A2 => n15131, B1 => n14899, B2 => 
                           n13671, ZN => n1781);
   U10956 : OAI22_X1 port map( A1 => n14909, A2 => n15062, B1 => n14908, B2 => 
                           n13812, ZN => n1790);
   U10957 : OAI22_X1 port map( A1 => n14909, A2 => n15065, B1 => n14908, B2 => 
                           n13813, ZN => n1791);
   U10958 : OAI22_X1 port map( A1 => n14909, A2 => n15068, B1 => n14908, B2 => 
                           n13814, ZN => n1792);
   U10959 : OAI22_X1 port map( A1 => n14909, A2 => n15071, B1 => n14908, B2 => 
                           n13815, ZN => n1793);
   U10960 : OAI22_X1 port map( A1 => n14909, A2 => n15074, B1 => n14908, B2 => 
                           n13816, ZN => n1794);
   U10961 : OAI22_X1 port map( A1 => n14910, A2 => n15077, B1 => n14908, B2 => 
                           n13817, ZN => n1795);
   U10962 : OAI22_X1 port map( A1 => n14910, A2 => n15080, B1 => n14908, B2 => 
                           n13818, ZN => n1796);
   U10963 : OAI22_X1 port map( A1 => n14910, A2 => n15083, B1 => n14908, B2 => 
                           n13819, ZN => n1797);
   U10964 : OAI22_X1 port map( A1 => n14910, A2 => n15086, B1 => n14908, B2 => 
                           n13820, ZN => n1798);
   U10965 : OAI22_X1 port map( A1 => n14910, A2 => n15089, B1 => n14908, B2 => 
                           n13821, ZN => n1799);
   U10966 : OAI22_X1 port map( A1 => n14911, A2 => n15092, B1 => n14908, B2 => 
                           n13822, ZN => n1800);
   U10967 : OAI22_X1 port map( A1 => n14911, A2 => n15095, B1 => n14908, B2 => 
                           n13823, ZN => n1801);
   U10968 : OAI22_X1 port map( A1 => n14911, A2 => n15098, B1 => n12007, B2 => 
                           n13712, ZN => n1802);
   U10969 : OAI22_X1 port map( A1 => n14911, A2 => n15101, B1 => n12007, B2 => 
                           n13713, ZN => n1803);
   U10970 : OAI22_X1 port map( A1 => n14911, A2 => n15104, B1 => n12007, B2 => 
                           n13714, ZN => n1804);
   U10971 : OAI22_X1 port map( A1 => n14912, A2 => n15107, B1 => n14908, B2 => 
                           n13715, ZN => n1805);
   U10972 : OAI22_X1 port map( A1 => n14912, A2 => n15110, B1 => n14908, B2 => 
                           n13716, ZN => n1806);
   U10973 : OAI22_X1 port map( A1 => n14912, A2 => n15113, B1 => n14908, B2 => 
                           n13717, ZN => n1807);
   U10974 : OAI22_X1 port map( A1 => n14912, A2 => n15116, B1 => n14908, B2 => 
                           n13718, ZN => n1808);
   U10975 : OAI22_X1 port map( A1 => n14912, A2 => n15119, B1 => n14908, B2 => 
                           n13719, ZN => n1809);
   U10976 : OAI22_X1 port map( A1 => n14913, A2 => n15122, B1 => n14908, B2 => 
                           n13720, ZN => n1810);
   U10977 : OAI22_X1 port map( A1 => n14913, A2 => n15125, B1 => n14908, B2 => 
                           n13721, ZN => n1811);
   U10978 : OAI22_X1 port map( A1 => n14913, A2 => n15128, B1 => n14908, B2 => 
                           n13722, ZN => n1812);
   U10979 : OAI22_X1 port map( A1 => n14913, A2 => n15131, B1 => n14908, B2 => 
                           n13723, ZN => n1813);
   U10980 : OAI22_X1 port map( A1 => n14918, A2 => n15062, B1 => n14917, B2 => 
                           n14142, ZN => n1822);
   U10981 : OAI22_X1 port map( A1 => n14918, A2 => n15065, B1 => n14917, B2 => 
                           n14143, ZN => n1823);
   U10982 : OAI22_X1 port map( A1 => n14918, A2 => n15068, B1 => n14917, B2 => 
                           n14144, ZN => n1824);
   U10983 : OAI22_X1 port map( A1 => n14918, A2 => n15071, B1 => n14917, B2 => 
                           n14145, ZN => n1825);
   U10984 : OAI22_X1 port map( A1 => n14918, A2 => n15074, B1 => n14917, B2 => 
                           n14146, ZN => n1826);
   U10985 : OAI22_X1 port map( A1 => n14919, A2 => n15077, B1 => n14917, B2 => 
                           n14147, ZN => n1827);
   U10986 : OAI22_X1 port map( A1 => n14919, A2 => n15080, B1 => n14917, B2 => 
                           n14148, ZN => n1828);
   U10987 : OAI22_X1 port map( A1 => n14919, A2 => n15083, B1 => n14917, B2 => 
                           n14149, ZN => n1829);
   U10988 : OAI22_X1 port map( A1 => n14919, A2 => n15086, B1 => n14917, B2 => 
                           n14150, ZN => n1830);
   U10989 : OAI22_X1 port map( A1 => n14919, A2 => n15089, B1 => n14917, B2 => 
                           n14151, ZN => n1831);
   U10990 : OAI22_X1 port map( A1 => n14920, A2 => n15092, B1 => n14917, B2 => 
                           n14152, ZN => n1832);
   U10991 : OAI22_X1 port map( A1 => n14920, A2 => n15095, B1 => n14917, B2 => 
                           n14153, ZN => n1833);
   U10992 : OAI22_X1 port map( A1 => n14920, A2 => n15098, B1 => n12005, B2 => 
                           n14154, ZN => n1834);
   U10993 : OAI22_X1 port map( A1 => n14920, A2 => n15101, B1 => n12005, B2 => 
                           n14155, ZN => n1835);
   U10994 : OAI22_X1 port map( A1 => n14920, A2 => n15104, B1 => n12005, B2 => 
                           n14156, ZN => n1836);
   U10995 : OAI22_X1 port map( A1 => n14921, A2 => n15107, B1 => n14917, B2 => 
                           n14157, ZN => n1837);
   U10996 : OAI22_X1 port map( A1 => n14921, A2 => n15110, B1 => n14917, B2 => 
                           n14158, ZN => n1838);
   U10997 : OAI22_X1 port map( A1 => n14921, A2 => n15113, B1 => n14917, B2 => 
                           n14159, ZN => n1839);
   U10998 : OAI22_X1 port map( A1 => n14921, A2 => n15116, B1 => n14917, B2 => 
                           n14160, ZN => n1840);
   U10999 : OAI22_X1 port map( A1 => n14921, A2 => n15119, B1 => n14917, B2 => 
                           n14161, ZN => n1841);
   U11000 : OAI22_X1 port map( A1 => n14922, A2 => n15122, B1 => n14917, B2 => 
                           n14162, ZN => n1842);
   U11001 : OAI22_X1 port map( A1 => n14922, A2 => n15125, B1 => n14917, B2 => 
                           n14163, ZN => n1843);
   U11002 : OAI22_X1 port map( A1 => n14922, A2 => n15128, B1 => n14917, B2 => 
                           n14164, ZN => n1844);
   U11003 : OAI22_X1 port map( A1 => n14922, A2 => n15131, B1 => n14917, B2 => 
                           n14165, ZN => n1845);
   U11004 : OAI22_X1 port map( A1 => n14972, A2 => n15061, B1 => n14971, B2 => 
                           n13740, ZN => n2014);
   U11005 : OAI22_X1 port map( A1 => n14972, A2 => n15064, B1 => n14971, B2 => 
                           n13741, ZN => n2015);
   U11006 : OAI22_X1 port map( A1 => n14972, A2 => n15067, B1 => n14971, B2 => 
                           n13742, ZN => n2016);
   U11007 : OAI22_X1 port map( A1 => n14972, A2 => n15070, B1 => n14971, B2 => 
                           n13743, ZN => n2017);
   U11008 : OAI22_X1 port map( A1 => n14972, A2 => n15073, B1 => n14971, B2 => 
                           n13744, ZN => n2018);
   U11009 : OAI22_X1 port map( A1 => n14973, A2 => n15076, B1 => n14971, B2 => 
                           n13745, ZN => n2019);
   U11010 : OAI22_X1 port map( A1 => n14973, A2 => n15079, B1 => n14971, B2 => 
                           n13746, ZN => n2020);
   U11011 : OAI22_X1 port map( A1 => n14973, A2 => n15082, B1 => n14971, B2 => 
                           n13747, ZN => n2021);
   U11012 : OAI22_X1 port map( A1 => n14973, A2 => n15085, B1 => n14971, B2 => 
                           n13748, ZN => n2022);
   U11013 : OAI22_X1 port map( A1 => n14973, A2 => n15088, B1 => n14971, B2 => 
                           n13749, ZN => n2023);
   U11014 : OAI22_X1 port map( A1 => n14974, A2 => n15091, B1 => n14971, B2 => 
                           n13750, ZN => n2024);
   U11015 : OAI22_X1 port map( A1 => n14974, A2 => n15094, B1 => n14971, B2 => 
                           n13751, ZN => n2025);
   U11016 : OAI22_X1 port map( A1 => n14974, A2 => n15097, B1 => n11998, B2 => 
                           n13672, ZN => n2026);
   U11017 : OAI22_X1 port map( A1 => n14974, A2 => n15100, B1 => n11998, B2 => 
                           n13673, ZN => n2027);
   U11018 : OAI22_X1 port map( A1 => n14974, A2 => n15103, B1 => n11998, B2 => 
                           n13674, ZN => n2028);
   U11019 : OAI22_X1 port map( A1 => n14975, A2 => n15106, B1 => n14971, B2 => 
                           n13675, ZN => n2029);
   U11020 : OAI22_X1 port map( A1 => n14975, A2 => n15109, B1 => n14971, B2 => 
                           n13676, ZN => n2030);
   U11021 : OAI22_X1 port map( A1 => n14975, A2 => n15112, B1 => n14971, B2 => 
                           n13677, ZN => n2031);
   U11022 : OAI22_X1 port map( A1 => n14975, A2 => n15115, B1 => n14971, B2 => 
                           n13678, ZN => n2032);
   U11023 : OAI22_X1 port map( A1 => n14975, A2 => n15118, B1 => n14971, B2 => 
                           n13679, ZN => n2033);
   U11024 : OAI22_X1 port map( A1 => n14976, A2 => n15121, B1 => n14971, B2 => 
                           n13680, ZN => n2034);
   U11025 : OAI22_X1 port map( A1 => n14976, A2 => n15124, B1 => n14971, B2 => 
                           n13681, ZN => n2035);
   U11026 : OAI22_X1 port map( A1 => n14976, A2 => n15127, B1 => n14971, B2 => 
                           n13682, ZN => n2036);
   U11027 : OAI22_X1 port map( A1 => n14976, A2 => n15130, B1 => n14971, B2 => 
                           n13683, ZN => n2037);
   U11028 : OAI22_X1 port map( A1 => n14981, A2 => n15061, B1 => n14980, B2 => 
                           n14094, ZN => n2046);
   U11029 : OAI22_X1 port map( A1 => n14981, A2 => n15064, B1 => n14980, B2 => 
                           n14095, ZN => n2047);
   U11030 : OAI22_X1 port map( A1 => n14981, A2 => n15067, B1 => n14980, B2 => 
                           n14096, ZN => n2048);
   U11031 : OAI22_X1 port map( A1 => n14981, A2 => n15070, B1 => n14980, B2 => 
                           n14097, ZN => n2049);
   U11032 : OAI22_X1 port map( A1 => n14981, A2 => n15073, B1 => n14980, B2 => 
                           n14098, ZN => n2050);
   U11033 : OAI22_X1 port map( A1 => n14982, A2 => n15076, B1 => n14980, B2 => 
                           n14099, ZN => n2051);
   U11034 : OAI22_X1 port map( A1 => n14982, A2 => n15079, B1 => n14980, B2 => 
                           n14100, ZN => n2052);
   U11035 : OAI22_X1 port map( A1 => n14982, A2 => n15082, B1 => n14980, B2 => 
                           n14101, ZN => n2053);
   U11036 : OAI22_X1 port map( A1 => n14982, A2 => n15085, B1 => n14980, B2 => 
                           n14102, ZN => n2054);
   U11037 : OAI22_X1 port map( A1 => n14982, A2 => n15088, B1 => n14980, B2 => 
                           n14103, ZN => n2055);
   U11038 : OAI22_X1 port map( A1 => n14983, A2 => n15091, B1 => n14980, B2 => 
                           n14104, ZN => n2056);
   U11039 : OAI22_X1 port map( A1 => n14983, A2 => n15094, B1 => n14980, B2 => 
                           n14105, ZN => n2057);
   U11040 : OAI22_X1 port map( A1 => n14983, A2 => n15097, B1 => n11997, B2 => 
                           n14106, ZN => n2058);
   U11041 : OAI22_X1 port map( A1 => n14983, A2 => n15100, B1 => n11997, B2 => 
                           n14107, ZN => n2059);
   U11042 : OAI22_X1 port map( A1 => n14983, A2 => n15103, B1 => n11997, B2 => 
                           n14108, ZN => n2060);
   U11043 : OAI22_X1 port map( A1 => n14984, A2 => n15106, B1 => n14980, B2 => 
                           n14109, ZN => n2061);
   U11044 : OAI22_X1 port map( A1 => n14984, A2 => n15109, B1 => n14980, B2 => 
                           n14110, ZN => n2062);
   U11045 : OAI22_X1 port map( A1 => n14984, A2 => n15112, B1 => n14980, B2 => 
                           n14111, ZN => n2063);
   U11046 : OAI22_X1 port map( A1 => n14984, A2 => n15115, B1 => n14980, B2 => 
                           n14112, ZN => n2064);
   U11047 : OAI22_X1 port map( A1 => n14984, A2 => n15118, B1 => n14980, B2 => 
                           n14113, ZN => n2065);
   U11048 : OAI22_X1 port map( A1 => n14985, A2 => n15121, B1 => n14980, B2 => 
                           n14114, ZN => n2066);
   U11049 : OAI22_X1 port map( A1 => n14985, A2 => n15124, B1 => n14980, B2 => 
                           n14115, ZN => n2067);
   U11050 : OAI22_X1 port map( A1 => n14985, A2 => n15127, B1 => n14980, B2 => 
                           n14116, ZN => n2068);
   U11051 : OAI22_X1 port map( A1 => n14985, A2 => n15130, B1 => n14980, B2 => 
                           n14117, ZN => n2069);
   U11052 : OAI22_X1 port map( A1 => n14990, A2 => n15061, B1 => n14989, B2 => 
                           n13832, ZN => n2078);
   U11053 : OAI22_X1 port map( A1 => n14990, A2 => n15064, B1 => n14989, B2 => 
                           n13833, ZN => n2079);
   U11054 : OAI22_X1 port map( A1 => n14990, A2 => n15067, B1 => n14989, B2 => 
                           n13834, ZN => n2080);
   U11055 : OAI22_X1 port map( A1 => n14990, A2 => n15070, B1 => n14989, B2 => 
                           n13835, ZN => n2081);
   U11056 : OAI22_X1 port map( A1 => n14990, A2 => n15073, B1 => n14989, B2 => 
                           n13836, ZN => n2082);
   U11057 : OAI22_X1 port map( A1 => n14991, A2 => n15076, B1 => n14989, B2 => 
                           n13837, ZN => n2083);
   U11058 : OAI22_X1 port map( A1 => n14991, A2 => n15079, B1 => n14989, B2 => 
                           n13838, ZN => n2084);
   U11059 : OAI22_X1 port map( A1 => n14991, A2 => n15082, B1 => n14989, B2 => 
                           n13839, ZN => n2085);
   U11060 : OAI22_X1 port map( A1 => n14991, A2 => n15085, B1 => n14989, B2 => 
                           n13840, ZN => n2086);
   U11061 : OAI22_X1 port map( A1 => n14991, A2 => n15088, B1 => n14989, B2 => 
                           n13841, ZN => n2087);
   U11062 : OAI22_X1 port map( A1 => n14992, A2 => n15091, B1 => n14989, B2 => 
                           n13842, ZN => n2088);
   U11063 : OAI22_X1 port map( A1 => n14992, A2 => n15094, B1 => n14989, B2 => 
                           n13843, ZN => n2089);
   U11064 : OAI22_X1 port map( A1 => n14992, A2 => n15097, B1 => n11995, B2 => 
                           n13768, ZN => n2090);
   U11065 : OAI22_X1 port map( A1 => n14992, A2 => n15100, B1 => n11995, B2 => 
                           n13769, ZN => n2091);
   U11066 : OAI22_X1 port map( A1 => n14992, A2 => n15103, B1 => n11995, B2 => 
                           n13770, ZN => n2092);
   U11067 : OAI22_X1 port map( A1 => n14993, A2 => n15106, B1 => n14989, B2 => 
                           n13771, ZN => n2093);
   U11068 : OAI22_X1 port map( A1 => n14993, A2 => n15109, B1 => n14989, B2 => 
                           n13772, ZN => n2094);
   U11069 : OAI22_X1 port map( A1 => n14993, A2 => n15112, B1 => n14989, B2 => 
                           n13773, ZN => n2095);
   U11070 : OAI22_X1 port map( A1 => n14993, A2 => n15115, B1 => n14989, B2 => 
                           n13774, ZN => n2096);
   U11071 : OAI22_X1 port map( A1 => n14993, A2 => n15118, B1 => n14989, B2 => 
                           n13775, ZN => n2097);
   U11072 : OAI22_X1 port map( A1 => n14994, A2 => n15121, B1 => n14989, B2 => 
                           n13776, ZN => n2098);
   U11073 : OAI22_X1 port map( A1 => n14994, A2 => n15124, B1 => n14989, B2 => 
                           n13777, ZN => n2099);
   U11074 : OAI22_X1 port map( A1 => n14994, A2 => n15127, B1 => n14989, B2 => 
                           n13778, ZN => n2100);
   U11075 : OAI22_X1 port map( A1 => n14994, A2 => n15130, B1 => n14989, B2 => 
                           n13779, ZN => n2101);
   U11076 : OAI22_X1 port map( A1 => n15044, A2 => n15061, B1 => n15043, B2 => 
                           n14086, ZN => n2270);
   U11077 : OAI22_X1 port map( A1 => n15044, A2 => n15064, B1 => n15043, B2 => 
                           n14087, ZN => n2271);
   U11078 : OAI22_X1 port map( A1 => n15044, A2 => n15067, B1 => n15043, B2 => 
                           n14088, ZN => n2272);
   U11079 : OAI22_X1 port map( A1 => n15044, A2 => n15070, B1 => n15043, B2 => 
                           n14089, ZN => n2273);
   U11080 : OAI22_X1 port map( A1 => n15044, A2 => n15073, B1 => n15043, B2 => 
                           n14090, ZN => n2274);
   U11081 : OAI22_X1 port map( A1 => n15045, A2 => n15076, B1 => n15043, B2 => 
                           n14091, ZN => n2275);
   U11082 : OAI22_X1 port map( A1 => n15045, A2 => n15079, B1 => n15043, B2 => 
                           n14092, ZN => n2276);
   U11083 : OAI22_X1 port map( A1 => n15045, A2 => n15082, B1 => n15043, B2 => 
                           n14093, ZN => n2277);
   U11084 : OAI22_X1 port map( A1 => n15045, A2 => n15085, B1 => n15043, B2 => 
                           n14070, ZN => n2278);
   U11085 : OAI22_X1 port map( A1 => n15045, A2 => n15088, B1 => n15043, B2 => 
                           n14071, ZN => n2279);
   U11086 : OAI22_X1 port map( A1 => n15046, A2 => n15091, B1 => n15043, B2 => 
                           n14072, ZN => n2280);
   U11087 : OAI22_X1 port map( A1 => n15046, A2 => n15094, B1 => n15043, B2 => 
                           n14073, ZN => n2281);
   U11088 : OAI22_X1 port map( A1 => n15046, A2 => n15097, B1 => n11985, B2 => 
                           n14074, ZN => n2282);
   U11089 : OAI22_X1 port map( A1 => n15046, A2 => n15100, B1 => n11985, B2 => 
                           n14075, ZN => n2283);
   U11090 : OAI22_X1 port map( A1 => n15046, A2 => n15103, B1 => n11985, B2 => 
                           n14076, ZN => n2284);
   U11091 : OAI22_X1 port map( A1 => n15047, A2 => n15106, B1 => n15043, B2 => 
                           n14077, ZN => n2285);
   U11092 : OAI22_X1 port map( A1 => n15047, A2 => n15109, B1 => n15043, B2 => 
                           n14078, ZN => n2286);
   U11093 : OAI22_X1 port map( A1 => n15047, A2 => n15112, B1 => n15043, B2 => 
                           n14079, ZN => n2287);
   U11094 : OAI22_X1 port map( A1 => n15047, A2 => n15115, B1 => n15043, B2 => 
                           n14080, ZN => n2288);
   U11095 : OAI22_X1 port map( A1 => n15047, A2 => n15118, B1 => n15043, B2 => 
                           n14081, ZN => n2289);
   U11096 : OAI22_X1 port map( A1 => n15048, A2 => n15121, B1 => n15043, B2 => 
                           n14082, ZN => n2290);
   U11097 : OAI22_X1 port map( A1 => n15048, A2 => n15124, B1 => n15043, B2 => 
                           n14083, ZN => n2291);
   U11098 : OAI22_X1 port map( A1 => n15048, A2 => n15127, B1 => n15043, B2 => 
                           n14084, ZN => n2292);
   U11099 : OAI22_X1 port map( A1 => n15048, A2 => n15130, B1 => n15043, B2 => 
                           n14085, ZN => n2293);
   U11100 : OAI22_X1 port map( A1 => n15053, A2 => n15061, B1 => n15052, B2 => 
                           n14118, ZN => n2302);
   U11101 : OAI22_X1 port map( A1 => n15053, A2 => n15064, B1 => n15052, B2 => 
                           n14119, ZN => n2303);
   U11102 : OAI22_X1 port map( A1 => n15053, A2 => n15067, B1 => n15052, B2 => 
                           n14120, ZN => n2304);
   U11103 : OAI22_X1 port map( A1 => n15053, A2 => n15070, B1 => n15052, B2 => 
                           n14121, ZN => n2305);
   U11104 : OAI22_X1 port map( A1 => n15053, A2 => n15073, B1 => n15052, B2 => 
                           n14122, ZN => n2306);
   U11105 : OAI22_X1 port map( A1 => n15054, A2 => n15076, B1 => n15052, B2 => 
                           n14123, ZN => n2307);
   U11106 : OAI22_X1 port map( A1 => n15054, A2 => n15079, B1 => n15052, B2 => 
                           n14124, ZN => n2308);
   U11107 : OAI22_X1 port map( A1 => n15054, A2 => n15082, B1 => n15052, B2 => 
                           n14125, ZN => n2309);
   U11108 : OAI22_X1 port map( A1 => n15054, A2 => n15085, B1 => n15052, B2 => 
                           n14126, ZN => n2310);
   U11109 : OAI22_X1 port map( A1 => n15054, A2 => n15088, B1 => n15052, B2 => 
                           n14127, ZN => n2311);
   U11110 : OAI22_X1 port map( A1 => n15055, A2 => n15091, B1 => n15052, B2 => 
                           n14128, ZN => n2312);
   U11111 : OAI22_X1 port map( A1 => n15055, A2 => n15094, B1 => n15052, B2 => 
                           n14129, ZN => n2313);
   U11112 : OAI22_X1 port map( A1 => n15055, A2 => n15097, B1 => n11983, B2 => 
                           n14130, ZN => n2314);
   U11113 : OAI22_X1 port map( A1 => n15055, A2 => n15100, B1 => n11983, B2 => 
                           n14131, ZN => n2315);
   U11114 : OAI22_X1 port map( A1 => n15055, A2 => n15103, B1 => n11983, B2 => 
                           n14132, ZN => n2316);
   U11115 : OAI22_X1 port map( A1 => n15056, A2 => n15106, B1 => n15052, B2 => 
                           n14133, ZN => n2317);
   U11116 : OAI22_X1 port map( A1 => n15056, A2 => n15109, B1 => n15052, B2 => 
                           n14134, ZN => n2318);
   U11117 : OAI22_X1 port map( A1 => n15056, A2 => n15112, B1 => n15052, B2 => 
                           n14135, ZN => n2319);
   U11118 : OAI22_X1 port map( A1 => n15056, A2 => n15115, B1 => n15052, B2 => 
                           n14136, ZN => n2320);
   U11119 : OAI22_X1 port map( A1 => n15056, A2 => n15118, B1 => n15052, B2 => 
                           n14137, ZN => n2321);
   U11120 : OAI22_X1 port map( A1 => n15057, A2 => n15121, B1 => n15052, B2 => 
                           n14138, ZN => n2322);
   U11121 : OAI22_X1 port map( A1 => n15057, A2 => n15124, B1 => n15052, B2 => 
                           n14139, ZN => n2323);
   U11122 : OAI22_X1 port map( A1 => n15057, A2 => n15127, B1 => n15052, B2 => 
                           n14140, ZN => n2324);
   U11123 : OAI22_X1 port map( A1 => n15057, A2 => n15130, B1 => n15052, B2 => 
                           n14141, ZN => n2325);
   U11124 : OAI22_X1 port map( A1 => n15155, A2 => n15061, B1 => n15154, B2 => 
                           n13844, ZN => n2334);
   U11125 : OAI22_X1 port map( A1 => n15155, A2 => n15064, B1 => n15154, B2 => 
                           n13845, ZN => n2335);
   U11126 : OAI22_X1 port map( A1 => n15155, A2 => n15067, B1 => n15154, B2 => 
                           n13846, ZN => n2336);
   U11127 : OAI22_X1 port map( A1 => n15155, A2 => n15070, B1 => n15154, B2 => 
                           n13847, ZN => n2337);
   U11128 : OAI22_X1 port map( A1 => n15155, A2 => n15073, B1 => n15154, B2 => 
                           n13848, ZN => n2338);
   U11129 : OAI22_X1 port map( A1 => n15156, A2 => n15076, B1 => n15154, B2 => 
                           n13849, ZN => n2339);
   U11130 : OAI22_X1 port map( A1 => n15156, A2 => n15079, B1 => n15154, B2 => 
                           n13850, ZN => n2340);
   U11131 : OAI22_X1 port map( A1 => n15156, A2 => n15082, B1 => n15154, B2 => 
                           n13851, ZN => n2341);
   U11132 : OAI22_X1 port map( A1 => n15156, A2 => n15085, B1 => n15154, B2 => 
                           n13852, ZN => n2342);
   U11133 : OAI22_X1 port map( A1 => n15156, A2 => n15088, B1 => n15154, B2 => 
                           n13853, ZN => n2343);
   U11134 : OAI22_X1 port map( A1 => n15157, A2 => n15091, B1 => n15154, B2 => 
                           n13854, ZN => n2344);
   U11135 : OAI22_X1 port map( A1 => n15157, A2 => n15094, B1 => n15154, B2 => 
                           n13855, ZN => n2345);
   U11136 : OAI22_X1 port map( A1 => n15157, A2 => n15097, B1 => n11949, B2 => 
                           n13780, ZN => n2346);
   U11137 : OAI22_X1 port map( A1 => n15157, A2 => n15100, B1 => n11949, B2 => 
                           n13781, ZN => n2347);
   U11138 : OAI22_X1 port map( A1 => n15157, A2 => n15103, B1 => n11949, B2 => 
                           n13782, ZN => n2348);
   U11139 : OAI22_X1 port map( A1 => n15158, A2 => n15106, B1 => n15154, B2 => 
                           n13783, ZN => n2349);
   U11140 : OAI22_X1 port map( A1 => n15158, A2 => n15109, B1 => n15154, B2 => 
                           n13784, ZN => n2350);
   U11141 : OAI22_X1 port map( A1 => n15158, A2 => n15112, B1 => n15154, B2 => 
                           n13785, ZN => n2351);
   U11142 : OAI22_X1 port map( A1 => n15158, A2 => n15115, B1 => n15154, B2 => 
                           n13786, ZN => n2352);
   U11143 : OAI22_X1 port map( A1 => n15158, A2 => n15118, B1 => n15154, B2 => 
                           n13787, ZN => n2353);
   U11144 : OAI22_X1 port map( A1 => n15159, A2 => n15121, B1 => n15154, B2 => 
                           n13788, ZN => n2354);
   U11145 : OAI22_X1 port map( A1 => n15159, A2 => n15124, B1 => n15154, B2 => 
                           n13789, ZN => n2355);
   U11146 : OAI22_X1 port map( A1 => n15159, A2 => n15127, B1 => n15154, B2 => 
                           n13790, ZN => n2356);
   U11147 : OAI22_X1 port map( A1 => n15159, A2 => n15130, B1 => n15154, B2 => 
                           n13791, ZN => n2357);
   U11148 : OAI22_X1 port map( A1 => n12025, A2 => n13637, B1 => n14781, B2 => 
                           n15066, ZN => n1343);
   U11149 : OAI22_X1 port map( A1 => n14780, A2 => n13638, B1 => n14781, B2 => 
                           n15069, ZN => n1344);
   U11150 : OAI22_X1 port map( A1 => n12025, A2 => n13639, B1 => n14781, B2 => 
                           n15072, ZN => n1345);
   U11151 : OAI22_X1 port map( A1 => n14780, A2 => n13640, B1 => n14782, B2 => 
                           n15075, ZN => n1346);
   U11152 : OAI22_X1 port map( A1 => n12025, A2 => n13641, B1 => n14782, B2 => 
                           n15078, ZN => n1347);
   U11153 : OAI22_X1 port map( A1 => n14780, A2 => n13642, B1 => n14782, B2 => 
                           n15081, ZN => n1348);
   U11154 : OAI22_X1 port map( A1 => n12025, A2 => n13643, B1 => n14782, B2 => 
                           n15084, ZN => n1349);
   U11155 : OAI22_X1 port map( A1 => n12025, A2 => n13724, B1 => n14783, B2 => 
                           n15087, ZN => n1350);
   U11156 : OAI22_X1 port map( A1 => n14780, A2 => n13725, B1 => n14783, B2 => 
                           n15090, ZN => n1351);
   U11157 : OAI22_X1 port map( A1 => n14780, A2 => n13726, B1 => n14783, B2 => 
                           n15093, ZN => n1352);
   U11158 : OAI22_X1 port map( A1 => n14780, A2 => n13636, B1 => n14788, B2 => 
                           n15153, ZN => n1372);
   U11159 : OAI22_X1 port map( A1 => n14780, A2 => n13727, B1 => n14788, B2 => 
                           n15165, ZN => n1373);
   U11160 : INV_X1 port map( A => n14578, ZN => n14669);
   U11161 : INV_X1 port map( A => n14580, ZN => n14659);
   U11162 : INV_X1 port map( A => n14578, ZN => n14670);
   U11163 : INV_X1 port map( A => n14580, ZN => n14660);
   U11164 : INV_X1 port map( A => n14579, ZN => n14767);
   U11165 : INV_X1 port map( A => n14581, ZN => n14757);
   U11166 : INV_X1 port map( A => n14579, ZN => n14768);
   U11167 : INV_X1 port map( A => n14581, ZN => n14758);
   U11168 : INV_X1 port map( A => n14582, ZN => n14661);
   U11169 : INV_X1 port map( A => n14583, ZN => n14759);
   U11170 : NAND2_X1 port map( A1 => n10990, A2 => n10991, ZN => n11982);
   U11171 : BUF_X1 port map( A => n12624, Z => n14667);
   U11172 : BUF_X1 port map( A => n12629, Z => n14657);
   U11173 : BUF_X1 port map( A => n12624, Z => n14666);
   U11174 : BUF_X1 port map( A => n12629, Z => n14656);
   U11175 : BUF_X1 port map( A => n12043, Z => n14765);
   U11176 : BUF_X1 port map( A => n12048, Z => n14755);
   U11177 : BUF_X1 port map( A => n12043, Z => n14764);
   U11178 : BUF_X1 port map( A => n12048, Z => n14754);
   U11179 : BUF_X1 port map( A => n12625, Z => n14663);
   U11180 : BUF_X1 port map( A => n12044, Z => n14761);
   U11181 : BUF_X1 port map( A => n12630, Z => n14654);
   U11182 : BUF_X1 port map( A => n12625, Z => n14664);
   U11183 : BUF_X1 port map( A => n12630, Z => n14653);
   U11184 : BUF_X1 port map( A => n12049, Z => n14752);
   U11185 : BUF_X1 port map( A => n12044, Z => n14762);
   U11186 : BUF_X1 port map( A => n12049, Z => n14751);
   U11187 : BUF_X1 port map( A => n12624, Z => n14668);
   U11188 : BUF_X1 port map( A => n12043, Z => n14766);
   U11189 : AND3_X1 port map( A1 => n11007, A2 => n11006, A3 => n14678, ZN => 
                           n13182);
   U11190 : AND3_X1 port map( A1 => n10999, A2 => n10998, A3 => n14776, ZN => 
                           n12601);
   U11191 : BUF_X1 port map( A => n12625, Z => n14665);
   U11192 : BUF_X1 port map( A => n12044, Z => n14763);
   U11193 : BUF_X1 port map( A => n10986, Z => n15169);
   U11194 : BUF_X1 port map( A => n10986, Z => n15170);
   U11195 : BUF_X1 port map( A => n12629, Z => n14658);
   U11196 : BUF_X1 port map( A => n12048, Z => n14756);
   U11197 : BUF_X1 port map( A => n10986, Z => n15167);
   U11198 : BUF_X1 port map( A => n10986, Z => n15166);
   U11199 : BUF_X1 port map( A => n11980, Z => n15062);
   U11200 : BUF_X1 port map( A => n11979, Z => n15065);
   U11201 : BUF_X1 port map( A => n11978, Z => n15068);
   U11202 : BUF_X1 port map( A => n11977, Z => n15071);
   U11203 : BUF_X1 port map( A => n11976, Z => n15074);
   U11204 : BUF_X1 port map( A => n11975, Z => n15077);
   U11205 : BUF_X1 port map( A => n11974, Z => n15080);
   U11206 : BUF_X1 port map( A => n11973, Z => n15083);
   U11207 : BUF_X1 port map( A => n11972, Z => n15086);
   U11208 : BUF_X1 port map( A => n11971, Z => n15089);
   U11209 : BUF_X1 port map( A => n11970, Z => n15092);
   U11210 : BUF_X1 port map( A => n11969, Z => n15095);
   U11211 : BUF_X1 port map( A => n11968, Z => n15098);
   U11212 : BUF_X1 port map( A => n11967, Z => n15101);
   U11213 : BUF_X1 port map( A => n11966, Z => n15104);
   U11214 : BUF_X1 port map( A => n11965, Z => n15107);
   U11215 : BUF_X1 port map( A => n11964, Z => n15110);
   U11216 : BUF_X1 port map( A => n11963, Z => n15113);
   U11217 : BUF_X1 port map( A => n11962, Z => n15116);
   U11218 : BUF_X1 port map( A => n11961, Z => n15119);
   U11219 : BUF_X1 port map( A => n11960, Z => n15122);
   U11220 : BUF_X1 port map( A => n11959, Z => n15125);
   U11221 : BUF_X1 port map( A => n11958, Z => n15128);
   U11222 : BUF_X1 port map( A => n11957, Z => n15131);
   U11223 : BUF_X1 port map( A => n11956, Z => n15134);
   U11224 : BUF_X1 port map( A => n11955, Z => n15137);
   U11225 : BUF_X1 port map( A => n11954, Z => n15140);
   U11226 : BUF_X1 port map( A => n11953, Z => n15143);
   U11227 : BUF_X1 port map( A => n11952, Z => n15146);
   U11228 : BUF_X1 port map( A => n11951, Z => n15149);
   U11229 : BUF_X1 port map( A => n11950, Z => n15152);
   U11230 : BUF_X1 port map( A => n11948, Z => n15164);
   U11231 : BUF_X1 port map( A => n11980, Z => n15061);
   U11232 : BUF_X1 port map( A => n11979, Z => n15064);
   U11233 : BUF_X1 port map( A => n11978, Z => n15067);
   U11234 : BUF_X1 port map( A => n11977, Z => n15070);
   U11235 : BUF_X1 port map( A => n11976, Z => n15073);
   U11236 : BUF_X1 port map( A => n11975, Z => n15076);
   U11237 : BUF_X1 port map( A => n11974, Z => n15079);
   U11238 : BUF_X1 port map( A => n11973, Z => n15082);
   U11239 : BUF_X1 port map( A => n11972, Z => n15085);
   U11240 : BUF_X1 port map( A => n11971, Z => n15088);
   U11241 : BUF_X1 port map( A => n11970, Z => n15091);
   U11242 : BUF_X1 port map( A => n11969, Z => n15094);
   U11243 : BUF_X1 port map( A => n11968, Z => n15097);
   U11244 : BUF_X1 port map( A => n11967, Z => n15100);
   U11245 : BUF_X1 port map( A => n11966, Z => n15103);
   U11246 : BUF_X1 port map( A => n11965, Z => n15106);
   U11247 : BUF_X1 port map( A => n11964, Z => n15109);
   U11248 : BUF_X1 port map( A => n11963, Z => n15112);
   U11249 : BUF_X1 port map( A => n11962, Z => n15115);
   U11250 : BUF_X1 port map( A => n11961, Z => n15118);
   U11251 : BUF_X1 port map( A => n11960, Z => n15121);
   U11252 : BUF_X1 port map( A => n11959, Z => n15124);
   U11253 : BUF_X1 port map( A => n11958, Z => n15127);
   U11254 : BUF_X1 port map( A => n11957, Z => n15130);
   U11255 : BUF_X1 port map( A => n11956, Z => n15133);
   U11256 : BUF_X1 port map( A => n11955, Z => n15136);
   U11257 : BUF_X1 port map( A => n11954, Z => n15139);
   U11258 : BUF_X1 port map( A => n11953, Z => n15142);
   U11259 : BUF_X1 port map( A => n11952, Z => n15145);
   U11260 : BUF_X1 port map( A => n11951, Z => n15148);
   U11261 : BUF_X1 port map( A => n11950, Z => n15151);
   U11262 : BUF_X1 port map( A => n11948, Z => n15163);
   U11263 : BUF_X1 port map( A => n10986, Z => n15168);
   U11264 : BUF_X1 port map( A => n12630, Z => n14655);
   U11265 : BUF_X1 port map( A => n12049, Z => n14753);
   U11266 : BUF_X1 port map( A => n12616, Z => n14676);
   U11267 : BUF_X1 port map( A => n12616, Z => n14677);
   U11268 : BUF_X1 port map( A => n12035, Z => n14774);
   U11269 : BUF_X1 port map( A => n12035, Z => n14775);
   U11270 : BUF_X1 port map( A => n12620, Z => n14673);
   U11271 : BUF_X1 port map( A => n12620, Z => n14674);
   U11272 : BUF_X1 port map( A => n12039, Z => n14771);
   U11273 : BUF_X1 port map( A => n12039, Z => n14772);
   U11274 : BUF_X1 port map( A => n11980, Z => n15063);
   U11275 : BUF_X1 port map( A => n11979, Z => n15066);
   U11276 : BUF_X1 port map( A => n11978, Z => n15069);
   U11277 : BUF_X1 port map( A => n11977, Z => n15072);
   U11278 : BUF_X1 port map( A => n11976, Z => n15075);
   U11279 : BUF_X1 port map( A => n11975, Z => n15078);
   U11280 : BUF_X1 port map( A => n11974, Z => n15081);
   U11281 : BUF_X1 port map( A => n11973, Z => n15084);
   U11282 : BUF_X1 port map( A => n11972, Z => n15087);
   U11283 : BUF_X1 port map( A => n11971, Z => n15090);
   U11284 : BUF_X1 port map( A => n11970, Z => n15093);
   U11285 : BUF_X1 port map( A => n11969, Z => n15096);
   U11286 : BUF_X1 port map( A => n11968, Z => n15099);
   U11287 : BUF_X1 port map( A => n11967, Z => n15102);
   U11288 : BUF_X1 port map( A => n11966, Z => n15105);
   U11289 : BUF_X1 port map( A => n11965, Z => n15108);
   U11290 : BUF_X1 port map( A => n11964, Z => n15111);
   U11291 : BUF_X1 port map( A => n11963, Z => n15114);
   U11292 : BUF_X1 port map( A => n11962, Z => n15117);
   U11293 : BUF_X1 port map( A => n11961, Z => n15120);
   U11294 : BUF_X1 port map( A => n11960, Z => n15123);
   U11295 : BUF_X1 port map( A => n11959, Z => n15126);
   U11296 : BUF_X1 port map( A => n11958, Z => n15129);
   U11297 : BUF_X1 port map( A => n11957, Z => n15132);
   U11298 : BUF_X1 port map( A => n11956, Z => n15135);
   U11299 : BUF_X1 port map( A => n11955, Z => n15138);
   U11300 : BUF_X1 port map( A => n11954, Z => n15141);
   U11301 : BUF_X1 port map( A => n11953, Z => n15144);
   U11302 : BUF_X1 port map( A => n11952, Z => n15147);
   U11303 : BUF_X1 port map( A => n11951, Z => n15150);
   U11304 : BUF_X1 port map( A => n11950, Z => n15153);
   U11305 : BUF_X1 port map( A => n11948, Z => n15165);
   U11306 : BUF_X1 port map( A => n12620, Z => n14675);
   U11307 : BUF_X1 port map( A => n12039, Z => n14773);
   U11308 : BUF_X1 port map( A => n12616, Z => n14678);
   U11309 : BUF_X1 port map( A => n12035, Z => n14776);
   U11310 : NAND2_X1 port map( A1 => n14663, A2 => n13181, ZN => n12615);
   U11311 : NAND2_X1 port map( A1 => n14663, A2 => n13183, ZN => n12631);
   U11312 : NAND2_X1 port map( A1 => n14761, A2 => n12600, ZN => n12034);
   U11313 : NAND2_X1 port map( A1 => n14761, A2 => n12602, ZN => n12050);
   U11314 : NAND2_X1 port map( A1 => n14668, A2 => n13181, ZN => n12632);
   U11315 : NAND2_X1 port map( A1 => n14668, A2 => n13183, ZN => n12634);
   U11316 : NAND2_X1 port map( A1 => n14766, A2 => n12600, ZN => n12051);
   U11317 : NAND2_X1 port map( A1 => n14766, A2 => n12602, ZN => n12053);
   U11318 : NAND2_X1 port map( A1 => n13181, A2 => n14582, ZN => n12647);
   U11319 : NAND2_X1 port map( A1 => n12600, A2 => n14583, ZN => n12066);
   U11320 : NAND2_X1 port map( A1 => n14578, A2 => n13181, ZN => n12635);
   U11321 : NAND2_X1 port map( A1 => n14580, A2 => n13181, ZN => n12645);
   U11322 : NAND2_X1 port map( A1 => n14579, A2 => n12600, ZN => n12054);
   U11323 : NAND2_X1 port map( A1 => n14581, A2 => n12600, ZN => n12064);
   U11324 : NAND2_X1 port map( A1 => n14578, A2 => n13183, ZN => n12637);
   U11325 : NAND2_X1 port map( A1 => n14580, A2 => n13183, ZN => n12648);
   U11326 : NAND2_X1 port map( A1 => n14579, A2 => n12602, ZN => n12056);
   U11327 : NAND2_X1 port map( A1 => n14581, A2 => n12602, ZN => n12067);
   U11328 : NAND2_X1 port map( A1 => n14578, A2 => n13182, ZN => n12638);
   U11329 : NAND2_X1 port map( A1 => n14580, A2 => n13182, ZN => n12646);
   U11330 : NAND2_X1 port map( A1 => n14579, A2 => n12601, ZN => n12057);
   U11331 : NAND2_X1 port map( A1 => n14581, A2 => n12601, ZN => n12065);
   U11332 : AND2_X1 port map( A1 => n13182, A2 => n14582, ZN => n12651);
   U11333 : AND2_X1 port map( A1 => n12601, A2 => n14583, ZN => n12070);
   U11334 : AND2_X1 port map( A1 => n14658, A2 => n13183, ZN => n12642);
   U11335 : AND2_X1 port map( A1 => n14658, A2 => n13181, ZN => n12654);
   U11336 : AND2_X1 port map( A1 => n14756, A2 => n12602, ZN => n12061);
   U11337 : AND2_X1 port map( A1 => n14756, A2 => n12600, ZN => n12073);
   U11338 : AND2_X1 port map( A1 => n14655, A2 => n13183, ZN => n12652);
   U11339 : AND2_X1 port map( A1 => n14655, A2 => n13181, ZN => n12657);
   U11340 : AND2_X1 port map( A1 => n14753, A2 => n12602, ZN => n12071);
   U11341 : AND2_X1 port map( A1 => n14753, A2 => n12600, ZN => n12076);
   U11342 : AND2_X1 port map( A1 => n14044, A2 => n13181, ZN => n12641);
   U11343 : AND2_X1 port map( A1 => n14045, A2 => n12600, ZN => n12060);
   U11344 : AND2_X1 port map( A1 => n14582, A2 => n13183, ZN => n12650);
   U11345 : AND2_X1 port map( A1 => n14583, A2 => n12602, ZN => n12069);
   U11346 : AND2_X1 port map( A1 => n14044, A2 => n13183, ZN => n12655);
   U11347 : AND2_X1 port map( A1 => n14045, A2 => n12602, ZN => n12074);
   U11348 : BUF_X1 port map( A => n12025, Z => n14780);
   U11349 : OAI21_X1 port map( B1 => n11988, B2 => n12022, A => n15171, ZN => 
                           n12025);
   U11350 : INV_X1 port map( A => n11987, ZN => n15042);
   U11351 : OAI21_X1 port map( B1 => n11981, B2 => n11988, A => n15170, ZN => 
                           n11987);
   U11352 : INV_X1 port map( A => n11985, ZN => n15051);
   U11353 : OAI21_X1 port map( B1 => n11981, B2 => n11986, A => n15170, ZN => 
                           n11985);
   U11354 : INV_X1 port map( A => n11983, ZN => n15060);
   U11355 : OAI21_X1 port map( B1 => n11981, B2 => n11984, A => n15171, ZN => 
                           n11983);
   U11356 : INV_X1 port map( A => n12024, ZN => n14799);
   U11357 : OAI21_X1 port map( B1 => n11986, B2 => n12022, A => n15168, ZN => 
                           n12024);
   U11358 : INV_X1 port map( A => n12023, ZN => n14808);
   U11359 : OAI21_X1 port map( B1 => n11984, B2 => n12022, A => n15168, ZN => 
                           n12023);
   U11360 : INV_X1 port map( A => n12021, ZN => n14817);
   U11361 : OAI21_X1 port map( B1 => n11982, B2 => n12022, A => n15168, ZN => 
                           n12021);
   U11362 : INV_X1 port map( A => n12020, ZN => n14826);
   U11363 : OAI21_X1 port map( B1 => n11988, B2 => n12017, A => n15169, ZN => 
                           n12020);
   U11364 : INV_X1 port map( A => n12019, ZN => n14835);
   U11365 : OAI21_X1 port map( B1 => n11986, B2 => n12017, A => n15169, ZN => 
                           n12019);
   U11366 : INV_X1 port map( A => n12018, ZN => n14844);
   U11367 : OAI21_X1 port map( B1 => n11984, B2 => n12017, A => n15169, ZN => 
                           n12018);
   U11368 : INV_X1 port map( A => n12016, ZN => n14853);
   U11369 : OAI21_X1 port map( B1 => n11982, B2 => n12017, A => n15169, ZN => 
                           n12016);
   U11370 : INV_X1 port map( A => n12015, ZN => n14862);
   U11371 : OAI21_X1 port map( B1 => n11988, B2 => n12012, A => n15169, ZN => 
                           n12015);
   U11372 : INV_X1 port map( A => n12014, ZN => n14871);
   U11373 : OAI21_X1 port map( B1 => n11986, B2 => n12012, A => n15169, ZN => 
                           n12014);
   U11374 : INV_X1 port map( A => n12013, ZN => n14880);
   U11375 : OAI21_X1 port map( B1 => n11984, B2 => n12012, A => n15169, ZN => 
                           n12013);
   U11376 : INV_X1 port map( A => n12011, ZN => n14889);
   U11377 : OAI21_X1 port map( B1 => n11982, B2 => n12012, A => n15169, ZN => 
                           n12011);
   U11378 : INV_X1 port map( A => n12009, ZN => n14898);
   U11379 : OAI21_X1 port map( B1 => n11988, B2 => n12006, A => n15169, ZN => 
                           n12009);
   U11380 : INV_X1 port map( A => n12008, ZN => n14907);
   U11381 : OAI21_X1 port map( B1 => n11986, B2 => n12006, A => n15169, ZN => 
                           n12008);
   U11382 : INV_X1 port map( A => n12007, ZN => n14916);
   U11383 : OAI21_X1 port map( B1 => n11984, B2 => n12006, A => n15169, ZN => 
                           n12007);
   U11384 : INV_X1 port map( A => n12004, ZN => n14934);
   U11385 : OAI21_X1 port map( B1 => n11988, B2 => n12001, A => n15169, ZN => 
                           n12004);
   U11386 : INV_X1 port map( A => n12003, ZN => n14943);
   U11387 : OAI21_X1 port map( B1 => n11986, B2 => n12001, A => n15170, ZN => 
                           n12003);
   U11388 : INV_X1 port map( A => n12002, ZN => n14952);
   U11389 : OAI21_X1 port map( B1 => n11984, B2 => n12001, A => n15170, ZN => 
                           n12002);
   U11390 : INV_X1 port map( A => n12000, ZN => n14961);
   U11391 : OAI21_X1 port map( B1 => n11982, B2 => n12001, A => n15170, ZN => 
                           n12000);
   U11392 : INV_X1 port map( A => n11999, ZN => n14970);
   U11393 : OAI21_X1 port map( B1 => n11988, B2 => n11996, A => n15170, ZN => 
                           n11999);
   U11394 : INV_X1 port map( A => n11998, ZN => n14979);
   U11395 : OAI21_X1 port map( B1 => n11986, B2 => n11996, A => n15170, ZN => 
                           n11998);
   U11396 : INV_X1 port map( A => n11997, ZN => n14988);
   U11397 : OAI21_X1 port map( B1 => n11984, B2 => n11996, A => n15170, ZN => 
                           n11997);
   U11398 : INV_X1 port map( A => n11995, ZN => n14997);
   U11399 : OAI21_X1 port map( B1 => n11982, B2 => n11996, A => n15170, ZN => 
                           n11995);
   U11400 : INV_X1 port map( A => n11994, ZN => n15006);
   U11401 : OAI21_X1 port map( B1 => n11988, B2 => n11991, A => n15170, ZN => 
                           n11994);
   U11402 : INV_X1 port map( A => n11993, ZN => n15015);
   U11403 : OAI21_X1 port map( B1 => n11986, B2 => n11991, A => n15170, ZN => 
                           n11993);
   U11404 : INV_X1 port map( A => n11992, ZN => n15024);
   U11405 : OAI21_X1 port map( B1 => n11984, B2 => n11991, A => n15170, ZN => 
                           n11992);
   U11406 : INV_X1 port map( A => n11990, ZN => n15033);
   U11407 : OAI21_X1 port map( B1 => n11982, B2 => n11991, A => n15170, ZN => 
                           n11990);
   U11408 : OAI221_X1 port map( B1 => n14070, B2 => n14679, C1 => n13200, C2 =>
                           n14677, A => n13040, ZN => n13039);
   U11409 : OAI21_X1 port map( B1 => n13041, B2 => n13042, A => n14673, ZN => 
                           n13040);
   U11410 : OAI221_X1 port map( B1 => n13724, B2 => n14662, C1 => n13880, C2 =>
                           n14659, A => n13044, ZN => n13041);
   U11411 : OAI221_X1 port map( B1 => n9523, B2 => n14671, C1 => n14166, C2 => 
                           n14669, A => n13043, ZN => n13042);
   U11412 : OAI221_X1 port map( B1 => n14071, B2 => n14679, C1 => n13201, C2 =>
                           n14677, A => n13023, ZN => n13022);
   U11413 : OAI21_X1 port map( B1 => n13024, B2 => n13025, A => n14673, ZN => 
                           n13023);
   U11414 : OAI221_X1 port map( B1 => n13725, B2 => n14662, C1 => n13881, C2 =>
                           n14659, A => n13027, ZN => n13024);
   U11415 : OAI221_X1 port map( B1 => n9522, B2 => n14671, C1 => n14167, C2 => 
                           n14669, A => n13026, ZN => n13025);
   U11416 : OAI221_X1 port map( B1 => n14072, B2 => n14679, C1 => n13202, C2 =>
                           n14677, A => n13006, ZN => n13005);
   U11417 : OAI21_X1 port map( B1 => n13007, B2 => n13008, A => n14673, ZN => 
                           n13006);
   U11418 : OAI221_X1 port map( B1 => n13726, B2 => n14662, C1 => n13882, C2 =>
                           n14659, A => n13010, ZN => n13007);
   U11419 : OAI221_X1 port map( B1 => n9521, B2 => n14671, C1 => n14168, C2 => 
                           n14669, A => n13009, ZN => n13008);
   U11420 : OAI221_X1 port map( B1 => n14073, B2 => n14679, C1 => n13203, C2 =>
                           n14677, A => n12989, ZN => n12988);
   U11421 : OAI21_X1 port map( B1 => n12990, B2 => n12991, A => n14673, ZN => 
                           n12989);
   U11422 : OAI221_X1 port map( B1 => n9648, B2 => n14662, C1 => n13883, C2 => 
                           n14659, A => n12993, ZN => n12990);
   U11423 : OAI221_X1 port map( B1 => n9520, B2 => n14671, C1 => n14169, C2 => 
                           n14669, A => n12992, ZN => n12991);
   U11424 : OAI221_X1 port map( B1 => n14074, B2 => n14680, C1 => n13204, C2 =>
                           n14677, A => n12972, ZN => n12971);
   U11425 : OAI21_X1 port map( B1 => n12973, B2 => n12974, A => n14674, ZN => 
                           n12972);
   U11426 : OAI221_X1 port map( B1 => n9647, B2 => n14661, C1 => n14170, C2 => 
                           n14660, A => n12976, ZN => n12973);
   U11427 : OAI221_X1 port map( B1 => n9519, B2 => n14672, C1 => n14171, C2 => 
                           n14670, A => n12975, ZN => n12974);
   U11428 : OAI221_X1 port map( B1 => n14075, B2 => n14680, C1 => n13205, C2 =>
                           n14677, A => n12955, ZN => n12954);
   U11429 : OAI21_X1 port map( B1 => n12956, B2 => n12957, A => n14674, ZN => 
                           n12955);
   U11430 : OAI221_X1 port map( B1 => n9646, B2 => n14661, C1 => n14172, C2 => 
                           n14660, A => n12959, ZN => n12956);
   U11431 : OAI221_X1 port map( B1 => n9518, B2 => n14672, C1 => n14173, C2 => 
                           n14670, A => n12958, ZN => n12957);
   U11432 : OAI221_X1 port map( B1 => n14076, B2 => n14680, C1 => n13206, C2 =>
                           n14677, A => n12938, ZN => n12937);
   U11433 : OAI21_X1 port map( B1 => n12939, B2 => n12940, A => n14674, ZN => 
                           n12938);
   U11434 : OAI221_X1 port map( B1 => n9645, B2 => n14661, C1 => n14174, C2 => 
                           n14660, A => n12942, ZN => n12939);
   U11435 : OAI221_X1 port map( B1 => n9517, B2 => n14672, C1 => n14175, C2 => 
                           n14670, A => n12941, ZN => n12940);
   U11436 : OAI221_X1 port map( B1 => n14077, B2 => n14680, C1 => n13207, C2 =>
                           n14677, A => n12921, ZN => n12920);
   U11437 : OAI21_X1 port map( B1 => n12922, B2 => n12923, A => n14674, ZN => 
                           n12921);
   U11438 : OAI221_X1 port map( B1 => n9644, B2 => n14661, C1 => n14176, C2 => 
                           n14660, A => n12925, ZN => n12922);
   U11439 : OAI221_X1 port map( B1 => n9516, B2 => n14672, C1 => n14177, C2 => 
                           n14670, A => n12924, ZN => n12923);
   U11440 : OAI221_X1 port map( B1 => n14078, B2 => n14680, C1 => n13208, C2 =>
                           n14677, A => n12904, ZN => n12903);
   U11441 : OAI21_X1 port map( B1 => n12905, B2 => n12906, A => n14674, ZN => 
                           n12904);
   U11442 : OAI221_X1 port map( B1 => n9643, B2 => n14661, C1 => n14178, C2 => 
                           n14660, A => n12908, ZN => n12905);
   U11443 : OAI221_X1 port map( B1 => n9515, B2 => n14672, C1 => n14179, C2 => 
                           n14670, A => n12907, ZN => n12906);
   U11444 : OAI221_X1 port map( B1 => n14079, B2 => n14680, C1 => n13209, C2 =>
                           n14677, A => n12887, ZN => n12886);
   U11445 : OAI21_X1 port map( B1 => n12888, B2 => n12889, A => n14674, ZN => 
                           n12887);
   U11446 : OAI221_X1 port map( B1 => n9642, B2 => n14661, C1 => n14180, C2 => 
                           n14660, A => n12891, ZN => n12888);
   U11447 : OAI221_X1 port map( B1 => n9514, B2 => n14672, C1 => n14181, C2 => 
                           n14670, A => n12890, ZN => n12889);
   U11448 : OAI221_X1 port map( B1 => n14080, B2 => n14680, C1 => n13210, C2 =>
                           n14677, A => n12870, ZN => n12869);
   U11449 : OAI21_X1 port map( B1 => n12871, B2 => n12872, A => n14674, ZN => 
                           n12870);
   U11450 : OAI221_X1 port map( B1 => n9641, B2 => n14661, C1 => n14182, C2 => 
                           n14660, A => n12874, ZN => n12871);
   U11451 : OAI221_X1 port map( B1 => n9513, B2 => n14672, C1 => n14183, C2 => 
                           n14670, A => n12873, ZN => n12872);
   U11452 : OAI221_X1 port map( B1 => n14081, B2 => n14680, C1 => n13211, C2 =>
                           n14676, A => n12853, ZN => n12852);
   U11453 : OAI21_X1 port map( B1 => n12854, B2 => n12855, A => n14674, ZN => 
                           n12853);
   U11454 : OAI221_X1 port map( B1 => n9640, B2 => n14661, C1 => n14184, C2 => 
                           n14660, A => n12857, ZN => n12854);
   U11455 : OAI221_X1 port map( B1 => n9512, B2 => n14672, C1 => n14185, C2 => 
                           n14670, A => n12856, ZN => n12855);
   U11456 : OAI221_X1 port map( B1 => n14082, B2 => n14680, C1 => n13212, C2 =>
                           n14676, A => n12836, ZN => n12835);
   U11457 : OAI21_X1 port map( B1 => n12837, B2 => n12838, A => n14674, ZN => 
                           n12836);
   U11458 : OAI221_X1 port map( B1 => n9639, B2 => n14661, C1 => n14186, C2 => 
                           n14660, A => n12840, ZN => n12837);
   U11459 : OAI221_X1 port map( B1 => n9511, B2 => n14672, C1 => n14187, C2 => 
                           n14670, A => n12839, ZN => n12838);
   U11460 : OAI221_X1 port map( B1 => n14083, B2 => n14680, C1 => n13213, C2 =>
                           n14676, A => n12819, ZN => n12818);
   U11461 : OAI21_X1 port map( B1 => n12820, B2 => n12821, A => n14674, ZN => 
                           n12819);
   U11462 : OAI221_X1 port map( B1 => n9638, B2 => n14661, C1 => n14188, C2 => 
                           n14660, A => n12823, ZN => n12820);
   U11463 : OAI221_X1 port map( B1 => n9510, B2 => n14672, C1 => n14189, C2 => 
                           n14670, A => n12822, ZN => n12821);
   U11464 : OAI221_X1 port map( B1 => n14084, B2 => n14680, C1 => n13214, C2 =>
                           n14676, A => n12802, ZN => n12801);
   U11465 : OAI21_X1 port map( B1 => n12803, B2 => n12804, A => n14674, ZN => 
                           n12802);
   U11466 : OAI221_X1 port map( B1 => n9637, B2 => n14661, C1 => n14190, C2 => 
                           n14660, A => n12806, ZN => n12803);
   U11467 : OAI221_X1 port map( B1 => n9509, B2 => n14672, C1 => n14191, C2 => 
                           n14670, A => n12805, ZN => n12804);
   U11468 : OAI221_X1 port map( B1 => n14085, B2 => n14680, C1 => n13215, C2 =>
                           n14676, A => n12785, ZN => n12784);
   U11469 : OAI21_X1 port map( B1 => n12786, B2 => n12787, A => n14674, ZN => 
                           n12785);
   U11470 : OAI221_X1 port map( B1 => n9636, B2 => n14661, C1 => n14192, C2 => 
                           n14660, A => n12789, ZN => n12786);
   U11471 : OAI221_X1 port map( B1 => n9508, B2 => n14672, C1 => n14193, C2 => 
                           n14670, A => n12788, ZN => n12787);
   U11472 : OAI221_X1 port map( B1 => n14070, B2 => n14777, C1 => n13230, C2 =>
                           n14775, A => n12459, ZN => n12458);
   U11473 : OAI21_X1 port map( B1 => n12460, B2 => n12461, A => n14771, ZN => 
                           n12459);
   U11474 : OAI221_X1 port map( B1 => n13724, B2 => n14760, C1 => n13880, C2 =>
                           n14757, A => n12463, ZN => n12460);
   U11475 : OAI221_X1 port map( B1 => n9523, B2 => n14769, C1 => n14166, C2 => 
                           n14767, A => n12462, ZN => n12461);
   U11476 : OAI221_X1 port map( B1 => n14071, B2 => n14777, C1 => n13231, C2 =>
                           n14775, A => n12442, ZN => n12441);
   U11477 : OAI21_X1 port map( B1 => n12443, B2 => n12444, A => n14771, ZN => 
                           n12442);
   U11478 : OAI221_X1 port map( B1 => n13725, B2 => n14760, C1 => n13881, C2 =>
                           n14757, A => n12446, ZN => n12443);
   U11479 : OAI221_X1 port map( B1 => n9522, B2 => n14769, C1 => n14167, C2 => 
                           n14767, A => n12445, ZN => n12444);
   U11480 : OAI221_X1 port map( B1 => n14072, B2 => n14777, C1 => n13232, C2 =>
                           n14775, A => n12425, ZN => n12424);
   U11481 : OAI21_X1 port map( B1 => n12426, B2 => n12427, A => n14771, ZN => 
                           n12425);
   U11482 : OAI221_X1 port map( B1 => n13726, B2 => n14760, C1 => n13882, C2 =>
                           n14757, A => n12429, ZN => n12426);
   U11483 : OAI221_X1 port map( B1 => n9521, B2 => n14769, C1 => n14168, C2 => 
                           n14767, A => n12428, ZN => n12427);
   U11484 : OAI221_X1 port map( B1 => n14073, B2 => n14777, C1 => n13233, C2 =>
                           n14775, A => n12408, ZN => n12407);
   U11485 : OAI21_X1 port map( B1 => n12409, B2 => n12410, A => n14771, ZN => 
                           n12408);
   U11486 : OAI221_X1 port map( B1 => n9648, B2 => n14760, C1 => n13883, C2 => 
                           n14757, A => n12412, ZN => n12409);
   U11487 : OAI221_X1 port map( B1 => n9520, B2 => n14769, C1 => n14169, C2 => 
                           n14767, A => n12411, ZN => n12410);
   U11488 : OAI221_X1 port map( B1 => n14074, B2 => n14778, C1 => n13234, C2 =>
                           n14775, A => n12391, ZN => n12390);
   U11489 : OAI21_X1 port map( B1 => n12392, B2 => n12393, A => n14772, ZN => 
                           n12391);
   U11490 : OAI221_X1 port map( B1 => n9647, B2 => n14759, C1 => n14170, C2 => 
                           n14758, A => n12395, ZN => n12392);
   U11491 : OAI221_X1 port map( B1 => n9519, B2 => n14770, C1 => n14171, C2 => 
                           n14768, A => n12394, ZN => n12393);
   U11492 : OAI221_X1 port map( B1 => n14075, B2 => n14778, C1 => n13235, C2 =>
                           n14775, A => n12374, ZN => n12373);
   U11493 : OAI21_X1 port map( B1 => n12375, B2 => n12376, A => n14772, ZN => 
                           n12374);
   U11494 : OAI221_X1 port map( B1 => n9646, B2 => n14759, C1 => n14172, C2 => 
                           n14758, A => n12378, ZN => n12375);
   U11495 : OAI221_X1 port map( B1 => n9518, B2 => n14770, C1 => n14173, C2 => 
                           n14768, A => n12377, ZN => n12376);
   U11496 : OAI221_X1 port map( B1 => n14076, B2 => n14778, C1 => n13236, C2 =>
                           n14775, A => n12357, ZN => n12356);
   U11497 : OAI21_X1 port map( B1 => n12358, B2 => n12359, A => n14772, ZN => 
                           n12357);
   U11498 : OAI221_X1 port map( B1 => n9645, B2 => n14759, C1 => n14174, C2 => 
                           n14758, A => n12361, ZN => n12358);
   U11499 : OAI221_X1 port map( B1 => n9517, B2 => n14770, C1 => n14175, C2 => 
                           n14768, A => n12360, ZN => n12359);
   U11500 : OAI221_X1 port map( B1 => n14077, B2 => n14778, C1 => n13237, C2 =>
                           n14775, A => n12340, ZN => n12339);
   U11501 : OAI21_X1 port map( B1 => n12341, B2 => n12342, A => n14772, ZN => 
                           n12340);
   U11502 : OAI221_X1 port map( B1 => n9644, B2 => n14759, C1 => n14176, C2 => 
                           n14758, A => n12344, ZN => n12341);
   U11503 : OAI221_X1 port map( B1 => n9516, B2 => n14770, C1 => n14177, C2 => 
                           n14768, A => n12343, ZN => n12342);
   U11504 : OAI221_X1 port map( B1 => n14078, B2 => n14778, C1 => n13238, C2 =>
                           n14775, A => n12323, ZN => n12322);
   U11505 : OAI21_X1 port map( B1 => n12324, B2 => n12325, A => n14772, ZN => 
                           n12323);
   U11506 : OAI221_X1 port map( B1 => n9643, B2 => n14759, C1 => n14178, C2 => 
                           n14758, A => n12327, ZN => n12324);
   U11507 : OAI221_X1 port map( B1 => n9515, B2 => n14770, C1 => n14179, C2 => 
                           n14768, A => n12326, ZN => n12325);
   U11508 : OAI221_X1 port map( B1 => n14079, B2 => n14778, C1 => n13239, C2 =>
                           n14775, A => n12306, ZN => n12305);
   U11509 : OAI21_X1 port map( B1 => n12307, B2 => n12308, A => n14772, ZN => 
                           n12306);
   U11510 : OAI221_X1 port map( B1 => n9642, B2 => n14759, C1 => n14180, C2 => 
                           n14758, A => n12310, ZN => n12307);
   U11511 : OAI221_X1 port map( B1 => n9514, B2 => n14770, C1 => n14181, C2 => 
                           n14768, A => n12309, ZN => n12308);
   U11512 : OAI221_X1 port map( B1 => n14080, B2 => n14778, C1 => n13240, C2 =>
                           n14775, A => n12289, ZN => n12288);
   U11513 : OAI21_X1 port map( B1 => n12290, B2 => n12291, A => n14772, ZN => 
                           n12289);
   U11514 : OAI221_X1 port map( B1 => n9641, B2 => n14759, C1 => n14182, C2 => 
                           n14758, A => n12293, ZN => n12290);
   U11515 : OAI221_X1 port map( B1 => n9513, B2 => n14770, C1 => n14183, C2 => 
                           n14768, A => n12292, ZN => n12291);
   U11516 : OAI221_X1 port map( B1 => n14081, B2 => n14778, C1 => n13241, C2 =>
                           n14774, A => n12272, ZN => n12271);
   U11517 : OAI21_X1 port map( B1 => n12273, B2 => n12274, A => n14772, ZN => 
                           n12272);
   U11518 : OAI221_X1 port map( B1 => n9640, B2 => n14759, C1 => n14184, C2 => 
                           n14758, A => n12276, ZN => n12273);
   U11519 : OAI221_X1 port map( B1 => n9512, B2 => n14770, C1 => n14185, C2 => 
                           n14768, A => n12275, ZN => n12274);
   U11520 : OAI221_X1 port map( B1 => n14082, B2 => n14778, C1 => n13242, C2 =>
                           n14774, A => n12255, ZN => n12254);
   U11521 : OAI21_X1 port map( B1 => n12256, B2 => n12257, A => n14772, ZN => 
                           n12255);
   U11522 : OAI221_X1 port map( B1 => n9639, B2 => n14759, C1 => n14186, C2 => 
                           n14758, A => n12259, ZN => n12256);
   U11523 : OAI221_X1 port map( B1 => n9511, B2 => n14770, C1 => n14187, C2 => 
                           n14768, A => n12258, ZN => n12257);
   U11524 : OAI221_X1 port map( B1 => n14083, B2 => n14778, C1 => n13243, C2 =>
                           n14774, A => n12238, ZN => n12237);
   U11525 : OAI21_X1 port map( B1 => n12239, B2 => n12240, A => n14772, ZN => 
                           n12238);
   U11526 : OAI221_X1 port map( B1 => n9638, B2 => n14759, C1 => n14188, C2 => 
                           n14758, A => n12242, ZN => n12239);
   U11527 : OAI221_X1 port map( B1 => n9510, B2 => n14770, C1 => n14189, C2 => 
                           n14768, A => n12241, ZN => n12240);
   U11528 : OAI221_X1 port map( B1 => n14084, B2 => n14778, C1 => n13244, C2 =>
                           n14774, A => n12221, ZN => n12220);
   U11529 : OAI21_X1 port map( B1 => n12222, B2 => n12223, A => n14772, ZN => 
                           n12221);
   U11530 : OAI221_X1 port map( B1 => n9637, B2 => n14759, C1 => n14190, C2 => 
                           n14758, A => n12225, ZN => n12222);
   U11531 : OAI221_X1 port map( B1 => n9509, B2 => n14770, C1 => n14191, C2 => 
                           n14768, A => n12224, ZN => n12223);
   U11532 : OAI221_X1 port map( B1 => n14085, B2 => n14778, C1 => n13245, C2 =>
                           n14774, A => n12204, ZN => n12203);
   U11533 : OAI21_X1 port map( B1 => n12205, B2 => n12206, A => n14772, ZN => 
                           n12204);
   U11534 : OAI221_X1 port map( B1 => n9636, B2 => n14759, C1 => n14192, C2 => 
                           n14758, A => n12208, ZN => n12205);
   U11535 : OAI221_X1 port map( B1 => n9508, B2 => n14770, C1 => n14193, C2 => 
                           n14768, A => n12207, ZN => n12206);
   U11536 : OAI221_X1 port map( B1 => n9627, B2 => n14611, C1 => n14194, C2 => 
                           n14608, A => n13187, ZN => n13185);
   U11537 : AOI22_X1 port map( A1 => n14605, A2 => n13948, B1 => n14604, B2 => 
                           n14354, ZN => n13187);
   U11538 : OAI221_X1 port map( B1 => n9626, B2 => n14611, C1 => n14195, C2 => 
                           n14608, A => n13167, ZN => n13165);
   U11539 : AOI22_X1 port map( A1 => n14605, A2 => n13949, B1 => n14604, B2 => 
                           n14355, ZN => n13167);
   U11540 : OAI221_X1 port map( B1 => n9625, B2 => n14611, C1 => n14196, C2 => 
                           n14608, A => n13150, ZN => n13148);
   U11541 : AOI22_X1 port map( A1 => n14605, A2 => n13950, B1 => n14604, B2 => 
                           n14356, ZN => n13150);
   U11542 : OAI221_X1 port map( B1 => n9624, B2 => n14611, C1 => n14197, C2 => 
                           n14608, A => n13133, ZN => n13131);
   U11543 : AOI22_X1 port map( A1 => n14605, A2 => n13951, B1 => n14604, B2 => 
                           n14357, ZN => n13133);
   U11544 : OAI221_X1 port map( B1 => n9623, B2 => n14611, C1 => n14198, C2 => 
                           n14608, A => n13116, ZN => n13114);
   U11545 : AOI22_X1 port map( A1 => n14605, A2 => n13952, B1 => n14604, B2 => 
                           n14358, ZN => n13116);
   U11546 : OAI221_X1 port map( B1 => n9622, B2 => n14611, C1 => n14199, C2 => 
                           n14608, A => n13099, ZN => n13097);
   U11547 : AOI22_X1 port map( A1 => n14605, A2 => n13953, B1 => n14604, B2 => 
                           n14359, ZN => n13099);
   U11548 : OAI221_X1 port map( B1 => n9621, B2 => n14611, C1 => n14200, C2 => 
                           n14608, A => n13082, ZN => n13080);
   U11549 : AOI22_X1 port map( A1 => n14605, A2 => n13954, B1 => n14604, B2 => 
                           n14360, ZN => n13082);
   U11550 : OAI221_X1 port map( B1 => n9620, B2 => n14611, C1 => n14201, C2 => 
                           n14608, A => n13065, ZN => n13063);
   U11551 : AOI22_X1 port map( A1 => n14605, A2 => n13955, B1 => n14604, B2 => 
                           n14361, ZN => n13065);
   U11552 : OAI221_X1 port map( B1 => n9619, B2 => n14611, C1 => n14202, C2 => 
                           n14608, A => n13048, ZN => n13046);
   U11553 : AOI22_X1 port map( A1 => n14605, A2 => n13956, B1 => n14603, B2 => 
                           n14362, ZN => n13048);
   U11554 : OAI221_X1 port map( B1 => n9618, B2 => n14611, C1 => n14203, C2 => 
                           n14608, A => n13031, ZN => n13029);
   U11555 : AOI22_X1 port map( A1 => n14605, A2 => n13957, B1 => n14603, B2 => 
                           n14363, ZN => n13031);
   U11556 : OAI221_X1 port map( B1 => n9617, B2 => n14611, C1 => n14204, C2 => 
                           n14608, A => n13014, ZN => n13012);
   U11557 : AOI22_X1 port map( A1 => n14605, A2 => n13958, B1 => n14603, B2 => 
                           n14364, ZN => n13014);
   U11558 : OAI221_X1 port map( B1 => n9616, B2 => n14611, C1 => n14205, C2 => 
                           n14608, A => n12997, ZN => n12995);
   U11559 : AOI22_X1 port map( A1 => n14605, A2 => n13959, B1 => n14603, B2 => 
                           n14365, ZN => n12997);
   U11560 : OAI221_X1 port map( B1 => n9615, B2 => n14612, C1 => n14206, C2 => 
                           n14609, A => n12980, ZN => n12978);
   U11561 : AOI22_X1 port map( A1 => n14606, A2 => n13960, B1 => n14603, B2 => 
                           n14366, ZN => n12980);
   U11562 : OAI221_X1 port map( B1 => n9614, B2 => n14612, C1 => n14207, C2 => 
                           n14609, A => n12963, ZN => n12961);
   U11563 : AOI22_X1 port map( A1 => n14606, A2 => n13961, B1 => n14603, B2 => 
                           n14367, ZN => n12963);
   U11564 : OAI221_X1 port map( B1 => n9613, B2 => n14612, C1 => n14208, C2 => 
                           n14609, A => n12946, ZN => n12944);
   U11565 : AOI22_X1 port map( A1 => n14606, A2 => n13962, B1 => n14603, B2 => 
                           n14368, ZN => n12946);
   U11566 : OAI221_X1 port map( B1 => n9612, B2 => n14612, C1 => n14209, C2 => 
                           n14609, A => n12929, ZN => n12927);
   U11567 : AOI22_X1 port map( A1 => n14606, A2 => n13963, B1 => n14603, B2 => 
                           n14369, ZN => n12929);
   U11568 : OAI221_X1 port map( B1 => n9611, B2 => n14612, C1 => n14210, C2 => 
                           n14609, A => n12912, ZN => n12910);
   U11569 : AOI22_X1 port map( A1 => n14606, A2 => n13964, B1 => n14603, B2 => 
                           n14370, ZN => n12912);
   U11570 : OAI221_X1 port map( B1 => n9610, B2 => n14612, C1 => n14211, C2 => 
                           n14609, A => n12895, ZN => n12893);
   U11571 : AOI22_X1 port map( A1 => n14606, A2 => n13965, B1 => n14603, B2 => 
                           n14371, ZN => n12895);
   U11572 : OAI221_X1 port map( B1 => n9609, B2 => n14612, C1 => n14212, C2 => 
                           n14609, A => n12878, ZN => n12876);
   U11573 : AOI22_X1 port map( A1 => n14606, A2 => n13966, B1 => n14603, B2 => 
                           n14372, ZN => n12878);
   U11574 : OAI221_X1 port map( B1 => n9608, B2 => n14612, C1 => n14213, C2 => 
                           n14609, A => n12861, ZN => n12859);
   U11575 : AOI22_X1 port map( A1 => n14606, A2 => n13967, B1 => n14603, B2 => 
                           n14373, ZN => n12861);
   U11576 : OAI221_X1 port map( B1 => n9607, B2 => n14612, C1 => n14214, C2 => 
                           n14609, A => n12844, ZN => n12842);
   U11577 : AOI22_X1 port map( A1 => n14606, A2 => n13968, B1 => n14602, B2 => 
                           n14374, ZN => n12844);
   U11578 : OAI221_X1 port map( B1 => n9606, B2 => n14612, C1 => n14215, C2 => 
                           n14609, A => n12827, ZN => n12825);
   U11579 : AOI22_X1 port map( A1 => n14606, A2 => n13969, B1 => n14602, B2 => 
                           n14375, ZN => n12827);
   U11580 : OAI221_X1 port map( B1 => n9605, B2 => n14612, C1 => n14216, C2 => 
                           n14609, A => n12810, ZN => n12808);
   U11581 : AOI22_X1 port map( A1 => n14606, A2 => n13970, B1 => n14602, B2 => 
                           n14376, ZN => n12810);
   U11582 : OAI221_X1 port map( B1 => n9604, B2 => n14612, C1 => n14217, C2 => 
                           n14609, A => n12793, ZN => n12791);
   U11583 : AOI22_X1 port map( A1 => n14606, A2 => n13971, B1 => n14602, B2 => 
                           n14377, ZN => n12793);
   U11584 : OAI221_X1 port map( B1 => n9627, B2 => n14709, C1 => n14194, C2 => 
                           n14706, A => n12606, ZN => n12604);
   U11585 : AOI22_X1 port map( A1 => n14703, A2 => n13948, B1 => n14702, B2 => 
                           n14354, ZN => n12606);
   U11586 : OAI221_X1 port map( B1 => n9626, B2 => n14709, C1 => n14195, C2 => 
                           n14706, A => n12586, ZN => n12584);
   U11587 : AOI22_X1 port map( A1 => n14703, A2 => n13949, B1 => n14702, B2 => 
                           n14355, ZN => n12586);
   U11588 : OAI221_X1 port map( B1 => n9625, B2 => n14709, C1 => n14196, C2 => 
                           n14706, A => n12569, ZN => n12567);
   U11589 : AOI22_X1 port map( A1 => n14703, A2 => n13950, B1 => n14702, B2 => 
                           n14356, ZN => n12569);
   U11590 : OAI221_X1 port map( B1 => n9624, B2 => n14709, C1 => n14197, C2 => 
                           n14706, A => n12552, ZN => n12550);
   U11591 : AOI22_X1 port map( A1 => n14703, A2 => n13951, B1 => n14702, B2 => 
                           n14357, ZN => n12552);
   U11592 : OAI221_X1 port map( B1 => n9623, B2 => n14709, C1 => n14198, C2 => 
                           n14706, A => n12535, ZN => n12533);
   U11593 : AOI22_X1 port map( A1 => n14703, A2 => n13952, B1 => n14702, B2 => 
                           n14358, ZN => n12535);
   U11594 : OAI221_X1 port map( B1 => n9622, B2 => n14709, C1 => n14199, C2 => 
                           n14706, A => n12518, ZN => n12516);
   U11595 : AOI22_X1 port map( A1 => n14703, A2 => n13953, B1 => n14702, B2 => 
                           n14359, ZN => n12518);
   U11596 : OAI221_X1 port map( B1 => n9621, B2 => n14709, C1 => n14200, C2 => 
                           n14706, A => n12501, ZN => n12499);
   U11597 : AOI22_X1 port map( A1 => n14703, A2 => n13954, B1 => n14702, B2 => 
                           n14360, ZN => n12501);
   U11598 : OAI221_X1 port map( B1 => n9620, B2 => n14709, C1 => n14201, C2 => 
                           n14706, A => n12484, ZN => n12482);
   U11599 : AOI22_X1 port map( A1 => n14703, A2 => n13955, B1 => n14702, B2 => 
                           n14361, ZN => n12484);
   U11600 : OAI221_X1 port map( B1 => n9619, B2 => n14709, C1 => n14202, C2 => 
                           n14706, A => n12467, ZN => n12465);
   U11601 : AOI22_X1 port map( A1 => n14703, A2 => n13956, B1 => n14701, B2 => 
                           n14362, ZN => n12467);
   U11602 : OAI221_X1 port map( B1 => n9618, B2 => n14709, C1 => n14203, C2 => 
                           n14706, A => n12450, ZN => n12448);
   U11603 : AOI22_X1 port map( A1 => n14703, A2 => n13957, B1 => n14701, B2 => 
                           n14363, ZN => n12450);
   U11604 : OAI221_X1 port map( B1 => n9617, B2 => n14709, C1 => n14204, C2 => 
                           n14706, A => n12433, ZN => n12431);
   U11605 : AOI22_X1 port map( A1 => n14703, A2 => n13958, B1 => n14701, B2 => 
                           n14364, ZN => n12433);
   U11606 : OAI221_X1 port map( B1 => n9616, B2 => n14709, C1 => n14205, C2 => 
                           n14706, A => n12416, ZN => n12414);
   U11607 : AOI22_X1 port map( A1 => n14703, A2 => n13959, B1 => n14701, B2 => 
                           n14365, ZN => n12416);
   U11608 : OAI221_X1 port map( B1 => n9615, B2 => n14710, C1 => n14206, C2 => 
                           n14707, A => n12399, ZN => n12397);
   U11609 : AOI22_X1 port map( A1 => n14704, A2 => n13960, B1 => n14701, B2 => 
                           n14366, ZN => n12399);
   U11610 : OAI221_X1 port map( B1 => n9614, B2 => n14710, C1 => n14207, C2 => 
                           n14707, A => n12382, ZN => n12380);
   U11611 : AOI22_X1 port map( A1 => n14704, A2 => n13961, B1 => n14701, B2 => 
                           n14367, ZN => n12382);
   U11612 : OAI221_X1 port map( B1 => n9613, B2 => n14710, C1 => n14208, C2 => 
                           n14707, A => n12365, ZN => n12363);
   U11613 : AOI22_X1 port map( A1 => n14704, A2 => n13962, B1 => n14701, B2 => 
                           n14368, ZN => n12365);
   U11614 : OAI221_X1 port map( B1 => n9612, B2 => n14710, C1 => n14209, C2 => 
                           n14707, A => n12348, ZN => n12346);
   U11615 : AOI22_X1 port map( A1 => n14704, A2 => n13963, B1 => n14701, B2 => 
                           n14369, ZN => n12348);
   U11616 : OAI221_X1 port map( B1 => n9611, B2 => n14710, C1 => n14210, C2 => 
                           n14707, A => n12331, ZN => n12329);
   U11617 : AOI22_X1 port map( A1 => n14704, A2 => n13964, B1 => n14701, B2 => 
                           n14370, ZN => n12331);
   U11618 : OAI221_X1 port map( B1 => n9610, B2 => n14710, C1 => n14211, C2 => 
                           n14707, A => n12314, ZN => n12312);
   U11619 : AOI22_X1 port map( A1 => n14704, A2 => n13965, B1 => n14701, B2 => 
                           n14371, ZN => n12314);
   U11620 : OAI221_X1 port map( B1 => n9609, B2 => n14710, C1 => n14212, C2 => 
                           n14707, A => n12297, ZN => n12295);
   U11621 : AOI22_X1 port map( A1 => n14704, A2 => n13966, B1 => n14701, B2 => 
                           n14372, ZN => n12297);
   U11622 : OAI221_X1 port map( B1 => n9608, B2 => n14710, C1 => n14213, C2 => 
                           n14707, A => n12280, ZN => n12278);
   U11623 : AOI22_X1 port map( A1 => n14704, A2 => n13967, B1 => n14701, B2 => 
                           n14373, ZN => n12280);
   U11624 : OAI221_X1 port map( B1 => n9607, B2 => n14710, C1 => n14214, C2 => 
                           n14707, A => n12263, ZN => n12261);
   U11625 : AOI22_X1 port map( A1 => n14704, A2 => n13968, B1 => n14700, B2 => 
                           n14374, ZN => n12263);
   U11626 : OAI221_X1 port map( B1 => n9606, B2 => n14710, C1 => n14215, C2 => 
                           n14707, A => n12246, ZN => n12244);
   U11627 : AOI22_X1 port map( A1 => n14704, A2 => n13969, B1 => n14700, B2 => 
                           n14375, ZN => n12246);
   U11628 : OAI221_X1 port map( B1 => n9605, B2 => n14710, C1 => n14216, C2 => 
                           n14707, A => n12229, ZN => n12227);
   U11629 : AOI22_X1 port map( A1 => n14704, A2 => n13970, B1 => n14700, B2 => 
                           n14376, ZN => n12229);
   U11630 : OAI221_X1 port map( B1 => n9604, B2 => n14710, C1 => n14217, C2 => 
                           n14707, A => n12212, ZN => n12210);
   U11631 : AOI22_X1 port map( A1 => n14704, A2 => n13971, B1 => n14700, B2 => 
                           n14377, ZN => n12212);
   U11632 : OAI22_X1 port map( A1 => n14940, A2 => n15134, B1 => n12003, B2 => 
                           n14028, ZN => n1910);
   U11633 : OAI22_X1 port map( A1 => n14941, A2 => n15137, B1 => n12003, B2 => 
                           n14029, ZN => n1911);
   U11634 : OAI22_X1 port map( A1 => n14941, A2 => n15140, B1 => n12003, B2 => 
                           n14030, ZN => n1912);
   U11635 : OAI22_X1 port map( A1 => n14941, A2 => n15143, B1 => n12003, B2 => 
                           n14031, ZN => n1913);
   U11636 : OAI22_X1 port map( A1 => n14941, A2 => n15146, B1 => n12003, B2 => 
                           n14032, ZN => n1914);
   U11637 : OAI22_X1 port map( A1 => n14941, A2 => n15149, B1 => n12003, B2 => 
                           n14033, ZN => n1915);
   U11638 : OAI22_X1 port map( A1 => n14942, A2 => n15152, B1 => n12003, B2 => 
                           n14034, ZN => n1916);
   U11639 : OAI22_X1 port map( A1 => n14942, A2 => n15164, B1 => n12003, B2 => 
                           n14035, ZN => n1917);
   U11640 : OAI22_X1 port map( A1 => n14949, A2 => n15134, B1 => n12002, B2 => 
                           n13988, ZN => n1942);
   U11641 : OAI22_X1 port map( A1 => n14950, A2 => n15137, B1 => n12002, B2 => 
                           n13989, ZN => n1943);
   U11642 : OAI22_X1 port map( A1 => n14950, A2 => n15140, B1 => n12002, B2 => 
                           n13990, ZN => n1944);
   U11643 : OAI22_X1 port map( A1 => n14950, A2 => n15143, B1 => n12002, B2 => 
                           n13991, ZN => n1945);
   U11644 : OAI22_X1 port map( A1 => n14950, A2 => n15146, B1 => n12002, B2 => 
                           n13992, ZN => n1946);
   U11645 : OAI22_X1 port map( A1 => n14950, A2 => n15149, B1 => n12002, B2 => 
                           n13993, ZN => n1947);
   U11646 : OAI22_X1 port map( A1 => n14951, A2 => n15152, B1 => n12002, B2 => 
                           n13994, ZN => n1948);
   U11647 : OAI22_X1 port map( A1 => n14951, A2 => n15164, B1 => n12002, B2 => 
                           n13995, ZN => n1949);
   U11648 : OAI22_X1 port map( A1 => n14958, A2 => n15134, B1 => n12000, B2 => 
                           n14012, ZN => n1974);
   U11649 : OAI22_X1 port map( A1 => n14959, A2 => n15137, B1 => n12000, B2 => 
                           n14013, ZN => n1975);
   U11650 : OAI22_X1 port map( A1 => n14959, A2 => n15140, B1 => n12000, B2 => 
                           n14014, ZN => n1976);
   U11651 : OAI22_X1 port map( A1 => n14959, A2 => n15143, B1 => n12000, B2 => 
                           n14015, ZN => n1977);
   U11652 : OAI22_X1 port map( A1 => n14959, A2 => n15146, B1 => n12000, B2 => 
                           n14016, ZN => n1978);
   U11653 : OAI22_X1 port map( A1 => n14959, A2 => n15149, B1 => n12000, B2 => 
                           n14017, ZN => n1979);
   U11654 : OAI22_X1 port map( A1 => n14960, A2 => n15152, B1 => n12000, B2 => 
                           n14018, ZN => n1980);
   U11655 : OAI22_X1 port map( A1 => n14960, A2 => n15164, B1 => n12000, B2 => 
                           n14019, ZN => n1981);
   U11656 : OAI22_X1 port map( A1 => n15003, A2 => n15133, B1 => n11994, B2 => 
                           n13996, ZN => n2134);
   U11657 : OAI22_X1 port map( A1 => n15004, A2 => n15136, B1 => n11994, B2 => 
                           n13997, ZN => n2135);
   U11658 : OAI22_X1 port map( A1 => n15004, A2 => n15139, B1 => n11994, B2 => 
                           n13998, ZN => n2136);
   U11659 : OAI22_X1 port map( A1 => n15004, A2 => n15142, B1 => n11994, B2 => 
                           n13999, ZN => n2137);
   U11660 : OAI22_X1 port map( A1 => n15004, A2 => n15145, B1 => n11994, B2 => 
                           n14000, ZN => n2138);
   U11661 : OAI22_X1 port map( A1 => n15004, A2 => n15148, B1 => n11994, B2 => 
                           n14001, ZN => n2139);
   U11662 : OAI22_X1 port map( A1 => n15005, A2 => n15151, B1 => n11994, B2 => 
                           n14002, ZN => n2140);
   U11663 : OAI22_X1 port map( A1 => n15005, A2 => n15163, B1 => n11994, B2 => 
                           n14003, ZN => n2141);
   U11664 : OAI22_X1 port map( A1 => n15012, A2 => n15133, B1 => n11993, B2 => 
                           n14036, ZN => n2166);
   U11665 : OAI22_X1 port map( A1 => n15013, A2 => n15136, B1 => n11993, B2 => 
                           n14037, ZN => n2167);
   U11666 : OAI22_X1 port map( A1 => n15013, A2 => n15139, B1 => n11993, B2 => 
                           n14038, ZN => n2168);
   U11667 : OAI22_X1 port map( A1 => n15013, A2 => n15142, B1 => n11993, B2 => 
                           n14039, ZN => n2169);
   U11668 : OAI22_X1 port map( A1 => n15013, A2 => n15145, B1 => n11993, B2 => 
                           n14040, ZN => n2170);
   U11669 : OAI22_X1 port map( A1 => n15013, A2 => n15148, B1 => n11993, B2 => 
                           n14041, ZN => n2171);
   U11670 : OAI22_X1 port map( A1 => n15014, A2 => n15151, B1 => n11993, B2 => 
                           n14042, ZN => n2172);
   U11671 : OAI22_X1 port map( A1 => n15014, A2 => n15163, B1 => n11993, B2 => 
                           n14043, ZN => n2173);
   U11672 : OAI22_X1 port map( A1 => n15021, A2 => n15133, B1 => n11992, B2 => 
                           n13980, ZN => n2198);
   U11673 : OAI22_X1 port map( A1 => n15022, A2 => n15136, B1 => n11992, B2 => 
                           n13981, ZN => n2199);
   U11674 : OAI22_X1 port map( A1 => n15022, A2 => n15139, B1 => n11992, B2 => 
                           n13982, ZN => n2200);
   U11675 : OAI22_X1 port map( A1 => n15022, A2 => n15142, B1 => n11992, B2 => 
                           n13983, ZN => n2201);
   U11676 : OAI22_X1 port map( A1 => n15022, A2 => n15145, B1 => n11992, B2 => 
                           n13984, ZN => n2202);
   U11677 : OAI22_X1 port map( A1 => n15022, A2 => n15148, B1 => n11992, B2 => 
                           n13985, ZN => n2203);
   U11678 : OAI22_X1 port map( A1 => n15023, A2 => n15151, B1 => n11992, B2 => 
                           n13986, ZN => n2204);
   U11679 : OAI22_X1 port map( A1 => n15023, A2 => n15163, B1 => n11992, B2 => 
                           n13987, ZN => n2205);
   U11680 : OAI22_X1 port map( A1 => n15030, A2 => n15133, B1 => n11990, B2 => 
                           n14020, ZN => n2230);
   U11681 : OAI22_X1 port map( A1 => n15031, A2 => n15136, B1 => n11990, B2 => 
                           n14021, ZN => n2231);
   U11682 : OAI22_X1 port map( A1 => n15031, A2 => n15139, B1 => n11990, B2 => 
                           n14022, ZN => n2232);
   U11683 : OAI22_X1 port map( A1 => n15031, A2 => n15142, B1 => n11990, B2 => 
                           n14023, ZN => n2233);
   U11684 : OAI22_X1 port map( A1 => n15031, A2 => n15145, B1 => n11990, B2 => 
                           n14024, ZN => n2234);
   U11685 : OAI22_X1 port map( A1 => n15031, A2 => n15148, B1 => n11990, B2 => 
                           n14025, ZN => n2235);
   U11686 : OAI22_X1 port map( A1 => n15032, A2 => n15151, B1 => n11990, B2 => 
                           n14026, ZN => n2236);
   U11687 : OAI22_X1 port map( A1 => n15032, A2 => n15163, B1 => n11990, B2 => 
                           n14027, ZN => n2237);
   U11688 : OAI22_X1 port map( A1 => n15039, A2 => n15133, B1 => n11987, B2 => 
                           n14004, ZN => n2262);
   U11689 : OAI22_X1 port map( A1 => n15040, A2 => n15136, B1 => n11987, B2 => 
                           n14005, ZN => n2263);
   U11690 : OAI22_X1 port map( A1 => n15040, A2 => n15139, B1 => n11987, B2 => 
                           n14006, ZN => n2264);
   U11691 : OAI22_X1 port map( A1 => n15040, A2 => n15142, B1 => n11987, B2 => 
                           n14007, ZN => n2265);
   U11692 : OAI22_X1 port map( A1 => n15040, A2 => n15145, B1 => n11987, B2 => 
                           n14008, ZN => n2266);
   U11693 : OAI22_X1 port map( A1 => n15040, A2 => n15148, B1 => n11987, B2 => 
                           n14009, ZN => n2267);
   U11694 : OAI22_X1 port map( A1 => n15041, A2 => n15151, B1 => n11987, B2 => 
                           n14010, ZN => n2268);
   U11695 : OAI22_X1 port map( A1 => n15041, A2 => n15163, B1 => n11987, B2 => 
                           n14011, ZN => n2269);
   U11696 : OAI22_X1 port map( A1 => n14796, A2 => n15135, B1 => n9603, B2 => 
                           n12024, ZN => n1398);
   U11697 : OAI22_X1 port map( A1 => n14797, A2 => n15138, B1 => n9602, B2 => 
                           n12024, ZN => n1399);
   U11698 : OAI22_X1 port map( A1 => n14797, A2 => n15141, B1 => n9601, B2 => 
                           n12024, ZN => n1400);
   U11699 : OAI22_X1 port map( A1 => n14797, A2 => n15144, B1 => n9600, B2 => 
                           n12024, ZN => n1401);
   U11700 : OAI22_X1 port map( A1 => n14797, A2 => n15147, B1 => n9599, B2 => 
                           n12024, ZN => n1402);
   U11701 : OAI22_X1 port map( A1 => n14797, A2 => n15150, B1 => n9598, B2 => 
                           n12024, ZN => n1403);
   U11702 : OAI22_X1 port map( A1 => n14798, A2 => n15153, B1 => n9597, B2 => 
                           n12024, ZN => n1404);
   U11703 : OAI22_X1 port map( A1 => n14798, A2 => n15165, B1 => n9596, B2 => 
                           n12024, ZN => n1405);
   U11704 : OAI22_X1 port map( A1 => n14805, A2 => n15135, B1 => n9571, B2 => 
                           n12023, ZN => n1430);
   U11705 : OAI22_X1 port map( A1 => n14806, A2 => n15138, B1 => n9570, B2 => 
                           n12023, ZN => n1431);
   U11706 : OAI22_X1 port map( A1 => n14806, A2 => n15141, B1 => n9569, B2 => 
                           n12023, ZN => n1432);
   U11707 : OAI22_X1 port map( A1 => n14806, A2 => n15144, B1 => n9568, B2 => 
                           n12023, ZN => n1433);
   U11708 : OAI22_X1 port map( A1 => n14806, A2 => n15147, B1 => n9567, B2 => 
                           n12023, ZN => n1434);
   U11709 : OAI22_X1 port map( A1 => n14806, A2 => n15150, B1 => n9566, B2 => 
                           n12023, ZN => n1435);
   U11710 : OAI22_X1 port map( A1 => n14807, A2 => n15153, B1 => n9565, B2 => 
                           n12023, ZN => n1436);
   U11711 : OAI22_X1 port map( A1 => n14807, A2 => n15165, B1 => n9564, B2 => 
                           n12023, ZN => n1437);
   U11712 : OAI22_X1 port map( A1 => n14814, A2 => n15135, B1 => n9539, B2 => 
                           n12021, ZN => n1462);
   U11713 : OAI22_X1 port map( A1 => n14815, A2 => n15138, B1 => n9538, B2 => 
                           n12021, ZN => n1463);
   U11714 : OAI22_X1 port map( A1 => n14815, A2 => n15141, B1 => n9537, B2 => 
                           n12021, ZN => n1464);
   U11715 : OAI22_X1 port map( A1 => n14815, A2 => n15144, B1 => n9536, B2 => 
                           n12021, ZN => n1465);
   U11716 : OAI22_X1 port map( A1 => n14815, A2 => n15147, B1 => n9535, B2 => 
                           n12021, ZN => n1466);
   U11717 : OAI22_X1 port map( A1 => n14815, A2 => n15150, B1 => n9534, B2 => 
                           n12021, ZN => n1467);
   U11718 : OAI22_X1 port map( A1 => n14816, A2 => n15153, B1 => n9533, B2 => 
                           n12021, ZN => n1468);
   U11719 : OAI22_X1 port map( A1 => n14816, A2 => n15165, B1 => n9532, B2 => 
                           n12021, ZN => n1469);
   U11720 : OAI22_X1 port map( A1 => n14823, A2 => n15135, B1 => n9507, B2 => 
                           n12020, ZN => n1494);
   U11721 : OAI22_X1 port map( A1 => n14824, A2 => n15138, B1 => n9506, B2 => 
                           n12020, ZN => n1495);
   U11722 : OAI22_X1 port map( A1 => n14824, A2 => n15141, B1 => n9505, B2 => 
                           n12020, ZN => n1496);
   U11723 : OAI22_X1 port map( A1 => n14824, A2 => n15144, B1 => n9504, B2 => 
                           n12020, ZN => n1497);
   U11724 : OAI22_X1 port map( A1 => n14824, A2 => n15147, B1 => n9503, B2 => 
                           n12020, ZN => n1498);
   U11725 : OAI22_X1 port map( A1 => n14824, A2 => n15150, B1 => n9502, B2 => 
                           n12020, ZN => n1499);
   U11726 : OAI22_X1 port map( A1 => n14825, A2 => n15153, B1 => n9501, B2 => 
                           n12020, ZN => n1500);
   U11727 : OAI22_X1 port map( A1 => n14825, A2 => n15165, B1 => n9500, B2 => 
                           n12020, ZN => n1501);
   U11728 : OAI22_X1 port map( A1 => n14832, A2 => n15135, B1 => n9475, B2 => 
                           n12019, ZN => n1526);
   U11729 : OAI22_X1 port map( A1 => n14833, A2 => n15138, B1 => n9474, B2 => 
                           n12019, ZN => n1527);
   U11730 : OAI22_X1 port map( A1 => n14833, A2 => n15141, B1 => n9473, B2 => 
                           n12019, ZN => n1528);
   U11731 : OAI22_X1 port map( A1 => n14833, A2 => n15144, B1 => n9472, B2 => 
                           n12019, ZN => n1529);
   U11732 : OAI22_X1 port map( A1 => n14833, A2 => n15147, B1 => n9471, B2 => 
                           n12019, ZN => n1530);
   U11733 : OAI22_X1 port map( A1 => n14833, A2 => n15150, B1 => n9470, B2 => 
                           n12019, ZN => n1531);
   U11734 : OAI22_X1 port map( A1 => n14834, A2 => n15153, B1 => n9469, B2 => 
                           n12019, ZN => n1532);
   U11735 : OAI22_X1 port map( A1 => n14834, A2 => n15165, B1 => n9468, B2 => 
                           n12019, ZN => n1533);
   U11736 : OAI22_X1 port map( A1 => n14841, A2 => n15135, B1 => n9443, B2 => 
                           n12018, ZN => n1558);
   U11737 : OAI22_X1 port map( A1 => n14842, A2 => n15138, B1 => n9442, B2 => 
                           n12018, ZN => n1559);
   U11738 : OAI22_X1 port map( A1 => n14842, A2 => n15141, B1 => n9441, B2 => 
                           n12018, ZN => n1560);
   U11739 : OAI22_X1 port map( A1 => n14842, A2 => n15144, B1 => n9440, B2 => 
                           n12018, ZN => n1561);
   U11740 : OAI22_X1 port map( A1 => n14842, A2 => n15147, B1 => n9439, B2 => 
                           n12018, ZN => n1562);
   U11741 : OAI22_X1 port map( A1 => n14842, A2 => n15150, B1 => n9438, B2 => 
                           n12018, ZN => n1563);
   U11742 : OAI22_X1 port map( A1 => n14843, A2 => n15153, B1 => n9437, B2 => 
                           n12018, ZN => n1564);
   U11743 : OAI22_X1 port map( A1 => n14843, A2 => n15165, B1 => n9436, B2 => 
                           n12018, ZN => n1565);
   U11744 : OAI22_X1 port map( A1 => n14850, A2 => n15135, B1 => n9411, B2 => 
                           n12016, ZN => n1590);
   U11745 : OAI22_X1 port map( A1 => n14851, A2 => n15138, B1 => n9410, B2 => 
                           n12016, ZN => n1591);
   U11746 : OAI22_X1 port map( A1 => n14851, A2 => n15141, B1 => n9409, B2 => 
                           n12016, ZN => n1592);
   U11747 : OAI22_X1 port map( A1 => n14851, A2 => n15144, B1 => n9408, B2 => 
                           n12016, ZN => n1593);
   U11748 : OAI22_X1 port map( A1 => n14851, A2 => n15147, B1 => n9407, B2 => 
                           n12016, ZN => n1594);
   U11749 : OAI22_X1 port map( A1 => n14851, A2 => n15150, B1 => n9406, B2 => 
                           n12016, ZN => n1595);
   U11750 : OAI22_X1 port map( A1 => n14852, A2 => n15153, B1 => n9405, B2 => 
                           n12016, ZN => n1596);
   U11751 : OAI22_X1 port map( A1 => n14852, A2 => n15165, B1 => n9404, B2 => 
                           n12016, ZN => n1597);
   U11752 : OAI22_X1 port map( A1 => n14931, A2 => n15134, B1 => n9123, B2 => 
                           n12004, ZN => n1878);
   U11753 : OAI22_X1 port map( A1 => n14932, A2 => n15137, B1 => n9122, B2 => 
                           n12004, ZN => n1879);
   U11754 : OAI22_X1 port map( A1 => n14932, A2 => n15140, B1 => n9121, B2 => 
                           n12004, ZN => n1880);
   U11755 : OAI22_X1 port map( A1 => n14932, A2 => n15143, B1 => n9120, B2 => 
                           n12004, ZN => n1881);
   U11756 : OAI22_X1 port map( A1 => n14932, A2 => n15146, B1 => n9119, B2 => 
                           n12004, ZN => n1882);
   U11757 : OAI22_X1 port map( A1 => n14932, A2 => n15149, B1 => n9118, B2 => 
                           n12004, ZN => n1883);
   U11758 : OAI22_X1 port map( A1 => n14933, A2 => n15152, B1 => n9117, B2 => 
                           n12004, ZN => n1884);
   U11759 : OAI22_X1 port map( A1 => n14933, A2 => n15164, B1 => n9116, B2 => 
                           n12004, ZN => n1885);
   U11760 : OAI22_X1 port map( A1 => n14967, A2 => n15133, B1 => n8995, B2 => 
                           n11999, ZN => n2006);
   U11761 : OAI22_X1 port map( A1 => n14968, A2 => n15136, B1 => n8994, B2 => 
                           n11999, ZN => n2007);
   U11762 : OAI22_X1 port map( A1 => n14968, A2 => n15139, B1 => n8993, B2 => 
                           n11999, ZN => n2008);
   U11763 : OAI22_X1 port map( A1 => n14968, A2 => n15142, B1 => n8992, B2 => 
                           n11999, ZN => n2009);
   U11764 : OAI22_X1 port map( A1 => n14968, A2 => n15145, B1 => n8991, B2 => 
                           n11999, ZN => n2010);
   U11765 : OAI22_X1 port map( A1 => n14968, A2 => n15148, B1 => n8990, B2 => 
                           n11999, ZN => n2011);
   U11766 : OAI22_X1 port map( A1 => n14969, A2 => n15151, B1 => n8989, B2 => 
                           n11999, ZN => n2012);
   U11767 : OAI22_X1 port map( A1 => n14969, A2 => n15163, B1 => n8988, B2 => 
                           n11999, ZN => n2013);
   U11768 : AOI22_X1 port map( A1 => n14668, A2 => n14258, B1 => n14663, B2 => 
                           n9670, ZN => n13179);
   U11769 : AOI22_X1 port map( A1 => n14658, A2 => n14259, B1 => n14655, B2 => 
                           n9897, ZN => n13180);
   U11770 : AOI22_X1 port map( A1 => n14668, A2 => n14260, B1 => n14663, B2 => 
                           n9671, ZN => n13162);
   U11771 : AOI22_X1 port map( A1 => n14658, A2 => n14261, B1 => n14655, B2 => 
                           n9899, ZN => n13163);
   U11772 : AOI22_X1 port map( A1 => n14668, A2 => n14262, B1 => n14663, B2 => 
                           n9672, ZN => n13145);
   U11773 : AOI22_X1 port map( A1 => n14658, A2 => n14263, B1 => n14655, B2 => 
                           n9901, ZN => n13146);
   U11774 : AOI22_X1 port map( A1 => n14668, A2 => n14264, B1 => n14663, B2 => 
                           n9673, ZN => n13128);
   U11775 : AOI22_X1 port map( A1 => n14658, A2 => n14265, B1 => n14655, B2 => 
                           n9903, ZN => n13129);
   U11776 : AOI22_X1 port map( A1 => n14668, A2 => n14266, B1 => n14663, B2 => 
                           n9674, ZN => n13111);
   U11777 : AOI22_X1 port map( A1 => n14658, A2 => n14267, B1 => n14655, B2 => 
                           n9905, ZN => n13112);
   U11778 : AOI22_X1 port map( A1 => n14668, A2 => n14268, B1 => n14663, B2 => 
                           n9675, ZN => n13094);
   U11779 : AOI22_X1 port map( A1 => n14658, A2 => n14269, B1 => n14655, B2 => 
                           n9907, ZN => n13095);
   U11780 : AOI22_X1 port map( A1 => n14668, A2 => n14270, B1 => n14663, B2 => 
                           n9676, ZN => n13077);
   U11781 : AOI22_X1 port map( A1 => n14658, A2 => n14271, B1 => n14655, B2 => 
                           n9909, ZN => n13078);
   U11782 : AOI22_X1 port map( A1 => n14668, A2 => n14272, B1 => n14663, B2 => 
                           n9677, ZN => n13060);
   U11783 : AOI22_X1 port map( A1 => n14658, A2 => n14273, B1 => n14655, B2 => 
                           n9911, ZN => n13061);
   U11784 : AOI22_X1 port map( A1 => n14667, A2 => n14274, B1 => n14663, B2 => 
                           n9678, ZN => n13043);
   U11785 : AOI22_X1 port map( A1 => n14657, A2 => n14275, B1 => n14654, B2 => 
                           n9913, ZN => n13044);
   U11786 : AOI22_X1 port map( A1 => n14667, A2 => n14276, B1 => n14664, B2 => 
                           n9679, ZN => n13026);
   U11787 : AOI22_X1 port map( A1 => n14657, A2 => n14277, B1 => n14654, B2 => 
                           n9915, ZN => n13027);
   U11788 : AOI22_X1 port map( A1 => n14667, A2 => n14278, B1 => n14664, B2 => 
                           n9680, ZN => n13009);
   U11789 : AOI22_X1 port map( A1 => n14657, A2 => n14279, B1 => n14654, B2 => 
                           n9917, ZN => n13010);
   U11790 : AOI22_X1 port map( A1 => n14667, A2 => n14280, B1 => n14664, B2 => 
                           n9681, ZN => n12992);
   U11791 : AOI22_X1 port map( A1 => n14657, A2 => n14281, B1 => n14654, B2 => 
                           n9919, ZN => n12993);
   U11792 : AOI22_X1 port map( A1 => n14667, A2 => n14282, B1 => n14664, B2 => 
                           n9682, ZN => n12975);
   U11793 : AOI22_X1 port map( A1 => n14657, A2 => n14283, B1 => n14654, B2 => 
                           n9921, ZN => n12976);
   U11794 : AOI22_X1 port map( A1 => n14667, A2 => n14284, B1 => n14664, B2 => 
                           n9683, ZN => n12958);
   U11795 : AOI22_X1 port map( A1 => n14657, A2 => n14285, B1 => n14654, B2 => 
                           n9923, ZN => n12959);
   U11796 : AOI22_X1 port map( A1 => n14667, A2 => n14286, B1 => n14664, B2 => 
                           n9684, ZN => n12941);
   U11797 : AOI22_X1 port map( A1 => n14657, A2 => n14287, B1 => n14654, B2 => 
                           n9925, ZN => n12942);
   U11798 : AOI22_X1 port map( A1 => n14667, A2 => n14288, B1 => n14664, B2 => 
                           n9685, ZN => n12924);
   U11799 : AOI22_X1 port map( A1 => n14657, A2 => n14289, B1 => n14654, B2 => 
                           n9927, ZN => n12925);
   U11800 : AOI22_X1 port map( A1 => n14667, A2 => n14290, B1 => n14664, B2 => 
                           n9686, ZN => n12907);
   U11801 : AOI22_X1 port map( A1 => n14657, A2 => n14291, B1 => n14654, B2 => 
                           n9929, ZN => n12908);
   U11802 : AOI22_X1 port map( A1 => n14667, A2 => n14292, B1 => n14664, B2 => 
                           n9687, ZN => n12890);
   U11803 : AOI22_X1 port map( A1 => n14657, A2 => n14293, B1 => n14654, B2 => 
                           n9931, ZN => n12891);
   U11804 : AOI22_X1 port map( A1 => n14667, A2 => n14294, B1 => n14664, B2 => 
                           n9688, ZN => n12873);
   U11805 : AOI22_X1 port map( A1 => n14657, A2 => n14295, B1 => n14654, B2 => 
                           n9933, ZN => n12874);
   U11806 : AOI22_X1 port map( A1 => n14667, A2 => n14296, B1 => n14664, B2 => 
                           n9689, ZN => n12856);
   U11807 : AOI22_X1 port map( A1 => n14657, A2 => n14297, B1 => n14654, B2 => 
                           n9935, ZN => n12857);
   U11808 : AOI22_X1 port map( A1 => n14666, A2 => n14298, B1 => n14664, B2 => 
                           n9690, ZN => n12839);
   U11809 : AOI22_X1 port map( A1 => n14656, A2 => n14299, B1 => n14653, B2 => 
                           n9937, ZN => n12840);
   U11810 : AOI22_X1 port map( A1 => n14666, A2 => n14300, B1 => n14665, B2 => 
                           n9691, ZN => n12822);
   U11811 : AOI22_X1 port map( A1 => n14656, A2 => n14301, B1 => n14653, B2 => 
                           n9939, ZN => n12823);
   U11812 : AOI22_X1 port map( A1 => n14666, A2 => n14302, B1 => n14665, B2 => 
                           n9692, ZN => n12805);
   U11813 : AOI22_X1 port map( A1 => n14656, A2 => n14303, B1 => n14653, B2 => 
                           n9941, ZN => n12806);
   U11814 : AOI22_X1 port map( A1 => n14666, A2 => n14304, B1 => n14665, B2 => 
                           n9693, ZN => n12788);
   U11815 : AOI22_X1 port map( A1 => n14656, A2 => n14305, B1 => n14653, B2 => 
                           n9943, ZN => n12789);
   U11816 : AOI22_X1 port map( A1 => n14666, A2 => n14306, B1 => n14665, B2 => 
                           n9694, ZN => n12771);
   U11817 : AOI22_X1 port map( A1 => n14656, A2 => n14307, B1 => n14653, B2 => 
                           n9945, ZN => n12772);
   U11818 : AOI22_X1 port map( A1 => n14666, A2 => n14308, B1 => n14665, B2 => 
                           n9695, ZN => n12754);
   U11819 : AOI22_X1 port map( A1 => n14656, A2 => n14309, B1 => n14653, B2 => 
                           n9947, ZN => n12755);
   U11820 : AOI22_X1 port map( A1 => n14666, A2 => n14310, B1 => n14665, B2 => 
                           n9696, ZN => n12737);
   U11821 : AOI22_X1 port map( A1 => n14656, A2 => n14311, B1 => n14653, B2 => 
                           n9949, ZN => n12738);
   U11822 : AOI22_X1 port map( A1 => n14666, A2 => n14312, B1 => n14665, B2 => 
                           n9697, ZN => n12720);
   U11823 : AOI22_X1 port map( A1 => n14656, A2 => n14313, B1 => n14653, B2 => 
                           n9951, ZN => n12721);
   U11824 : AOI22_X1 port map( A1 => n14666, A2 => n14314, B1 => n14665, B2 => 
                           n9698, ZN => n12703);
   U11825 : AOI22_X1 port map( A1 => n14656, A2 => n14315, B1 => n14653, B2 => 
                           n9953, ZN => n12704);
   U11826 : AOI22_X1 port map( A1 => n14666, A2 => n14316, B1 => n14665, B2 => 
                           n9699, ZN => n12686);
   U11827 : AOI22_X1 port map( A1 => n14656, A2 => n14317, B1 => n14653, B2 => 
                           n9955, ZN => n12687);
   U11828 : AOI22_X1 port map( A1 => n14666, A2 => n14318, B1 => n14665, B2 => 
                           n9700, ZN => n12669);
   U11829 : AOI22_X1 port map( A1 => n14656, A2 => n14319, B1 => n14653, B2 => 
                           n9893, ZN => n12670);
   U11830 : AOI22_X1 port map( A1 => n14666, A2 => n14320, B1 => n14665, B2 => 
                           n9701, ZN => n12623);
   U11831 : AOI22_X1 port map( A1 => n14656, A2 => n14321, B1 => n14653, B2 => 
                           n9895, ZN => n12628);
   U11832 : AOI22_X1 port map( A1 => n14766, A2 => n14258, B1 => n14761, B2 => 
                           n9670, ZN => n12598);
   U11833 : AOI22_X1 port map( A1 => n14756, A2 => n14259, B1 => n14753, B2 => 
                           n9897, ZN => n12599);
   U11834 : AOI22_X1 port map( A1 => n14766, A2 => n14260, B1 => n14761, B2 => 
                           n9671, ZN => n12581);
   U11835 : AOI22_X1 port map( A1 => n14756, A2 => n14261, B1 => n14753, B2 => 
                           n9899, ZN => n12582);
   U11836 : AOI22_X1 port map( A1 => n14766, A2 => n14262, B1 => n14761, B2 => 
                           n9672, ZN => n12564);
   U11837 : AOI22_X1 port map( A1 => n14756, A2 => n14263, B1 => n14753, B2 => 
                           n9901, ZN => n12565);
   U11838 : AOI22_X1 port map( A1 => n14766, A2 => n14264, B1 => n14761, B2 => 
                           n9673, ZN => n12547);
   U11839 : AOI22_X1 port map( A1 => n14756, A2 => n14265, B1 => n14753, B2 => 
                           n9903, ZN => n12548);
   U11840 : AOI22_X1 port map( A1 => n14766, A2 => n14266, B1 => n14761, B2 => 
                           n9674, ZN => n12530);
   U11841 : AOI22_X1 port map( A1 => n14756, A2 => n14267, B1 => n14753, B2 => 
                           n9905, ZN => n12531);
   U11842 : AOI22_X1 port map( A1 => n14766, A2 => n14268, B1 => n14761, B2 => 
                           n9675, ZN => n12513);
   U11843 : AOI22_X1 port map( A1 => n14756, A2 => n14269, B1 => n14753, B2 => 
                           n9907, ZN => n12514);
   U11844 : AOI22_X1 port map( A1 => n14766, A2 => n14270, B1 => n14761, B2 => 
                           n9676, ZN => n12496);
   U11845 : AOI22_X1 port map( A1 => n14756, A2 => n14271, B1 => n14753, B2 => 
                           n9909, ZN => n12497);
   U11846 : AOI22_X1 port map( A1 => n14766, A2 => n14272, B1 => n14761, B2 => 
                           n9677, ZN => n12479);
   U11847 : AOI22_X1 port map( A1 => n14756, A2 => n14273, B1 => n14753, B2 => 
                           n9911, ZN => n12480);
   U11848 : AOI22_X1 port map( A1 => n14765, A2 => n14274, B1 => n14761, B2 => 
                           n9678, ZN => n12462);
   U11849 : AOI22_X1 port map( A1 => n14755, A2 => n14275, B1 => n14752, B2 => 
                           n9913, ZN => n12463);
   U11850 : AOI22_X1 port map( A1 => n14765, A2 => n14276, B1 => n14762, B2 => 
                           n9679, ZN => n12445);
   U11851 : AOI22_X1 port map( A1 => n14755, A2 => n14277, B1 => n14752, B2 => 
                           n9915, ZN => n12446);
   U11852 : AOI22_X1 port map( A1 => n14765, A2 => n14278, B1 => n14762, B2 => 
                           n9680, ZN => n12428);
   U11853 : AOI22_X1 port map( A1 => n14755, A2 => n14279, B1 => n14752, B2 => 
                           n9917, ZN => n12429);
   U11854 : AOI22_X1 port map( A1 => n14765, A2 => n14280, B1 => n14762, B2 => 
                           n9681, ZN => n12411);
   U11855 : AOI22_X1 port map( A1 => n14755, A2 => n14281, B1 => n14752, B2 => 
                           n9919, ZN => n12412);
   U11856 : AOI22_X1 port map( A1 => n14765, A2 => n14282, B1 => n14762, B2 => 
                           n9682, ZN => n12394);
   U11857 : AOI22_X1 port map( A1 => n14755, A2 => n14283, B1 => n14752, B2 => 
                           n9921, ZN => n12395);
   U11858 : AOI22_X1 port map( A1 => n14765, A2 => n14284, B1 => n14762, B2 => 
                           n9683, ZN => n12377);
   U11859 : AOI22_X1 port map( A1 => n14755, A2 => n14285, B1 => n14752, B2 => 
                           n9923, ZN => n12378);
   U11860 : AOI22_X1 port map( A1 => n14765, A2 => n14286, B1 => n14762, B2 => 
                           n9684, ZN => n12360);
   U11861 : AOI22_X1 port map( A1 => n14755, A2 => n14287, B1 => n14752, B2 => 
                           n9925, ZN => n12361);
   U11862 : AOI22_X1 port map( A1 => n14765, A2 => n14288, B1 => n14762, B2 => 
                           n9685, ZN => n12343);
   U11863 : AOI22_X1 port map( A1 => n14755, A2 => n14289, B1 => n14752, B2 => 
                           n9927, ZN => n12344);
   U11864 : AOI22_X1 port map( A1 => n14765, A2 => n14290, B1 => n14762, B2 => 
                           n9686, ZN => n12326);
   U11865 : AOI22_X1 port map( A1 => n14755, A2 => n14291, B1 => n14752, B2 => 
                           n9929, ZN => n12327);
   U11866 : AOI22_X1 port map( A1 => n14765, A2 => n14292, B1 => n14762, B2 => 
                           n9687, ZN => n12309);
   U11867 : AOI22_X1 port map( A1 => n14755, A2 => n14293, B1 => n14752, B2 => 
                           n9931, ZN => n12310);
   U11868 : AOI22_X1 port map( A1 => n14765, A2 => n14294, B1 => n14762, B2 => 
                           n9688, ZN => n12292);
   U11869 : AOI22_X1 port map( A1 => n14755, A2 => n14295, B1 => n14752, B2 => 
                           n9933, ZN => n12293);
   U11870 : AOI22_X1 port map( A1 => n14765, A2 => n14296, B1 => n14762, B2 => 
                           n9689, ZN => n12275);
   U11871 : AOI22_X1 port map( A1 => n14755, A2 => n14297, B1 => n14752, B2 => 
                           n9935, ZN => n12276);
   U11872 : AOI22_X1 port map( A1 => n14764, A2 => n14298, B1 => n14762, B2 => 
                           n9690, ZN => n12258);
   U11873 : AOI22_X1 port map( A1 => n14754, A2 => n14299, B1 => n14751, B2 => 
                           n9937, ZN => n12259);
   U11874 : AOI22_X1 port map( A1 => n14764, A2 => n14300, B1 => n14763, B2 => 
                           n9691, ZN => n12241);
   U11875 : AOI22_X1 port map( A1 => n14754, A2 => n14301, B1 => n14751, B2 => 
                           n9939, ZN => n12242);
   U11876 : AOI22_X1 port map( A1 => n14764, A2 => n14302, B1 => n14763, B2 => 
                           n9692, ZN => n12224);
   U11877 : AOI22_X1 port map( A1 => n14754, A2 => n14303, B1 => n14751, B2 => 
                           n9941, ZN => n12225);
   U11878 : AOI22_X1 port map( A1 => n14764, A2 => n14304, B1 => n14763, B2 => 
                           n9693, ZN => n12207);
   U11879 : AOI22_X1 port map( A1 => n14754, A2 => n14305, B1 => n14751, B2 => 
                           n9943, ZN => n12208);
   U11880 : AOI22_X1 port map( A1 => n14764, A2 => n14306, B1 => n14763, B2 => 
                           n9694, ZN => n12190);
   U11881 : AOI22_X1 port map( A1 => n14754, A2 => n14307, B1 => n14751, B2 => 
                           n9945, ZN => n12191);
   U11882 : AOI22_X1 port map( A1 => n14764, A2 => n14308, B1 => n14763, B2 => 
                           n9695, ZN => n12173);
   U11883 : AOI22_X1 port map( A1 => n14754, A2 => n14309, B1 => n14751, B2 => 
                           n9947, ZN => n12174);
   U11884 : AOI22_X1 port map( A1 => n14764, A2 => n14310, B1 => n14763, B2 => 
                           n9696, ZN => n12156);
   U11885 : AOI22_X1 port map( A1 => n14754, A2 => n14311, B1 => n14751, B2 => 
                           n9949, ZN => n12157);
   U11886 : AOI22_X1 port map( A1 => n14764, A2 => n14312, B1 => n14763, B2 => 
                           n9697, ZN => n12139);
   U11887 : AOI22_X1 port map( A1 => n14754, A2 => n14313, B1 => n14751, B2 => 
                           n9951, ZN => n12140);
   U11888 : AOI22_X1 port map( A1 => n14764, A2 => n14314, B1 => n14763, B2 => 
                           n9698, ZN => n12122);
   U11889 : AOI22_X1 port map( A1 => n14754, A2 => n14315, B1 => n14751, B2 => 
                           n9953, ZN => n12123);
   U11890 : AOI22_X1 port map( A1 => n14764, A2 => n14316, B1 => n14763, B2 => 
                           n9699, ZN => n12105);
   U11891 : AOI22_X1 port map( A1 => n14754, A2 => n14317, B1 => n14751, B2 => 
                           n9955, ZN => n12106);
   U11892 : AOI22_X1 port map( A1 => n14764, A2 => n14318, B1 => n14763, B2 => 
                           n9700, ZN => n12088);
   U11893 : AOI22_X1 port map( A1 => n14754, A2 => n14319, B1 => n14751, B2 => 
                           n9893, ZN => n12089);
   U11894 : AOI22_X1 port map( A1 => n14764, A2 => n14320, B1 => n14763, B2 => 
                           n9701, ZN => n12042);
   U11895 : AOI22_X1 port map( A1 => n14754, A2 => n14321, B1 => n14751, B2 => 
                           n9895, ZN => n12047);
   U11896 : OAI221_X1 port map( B1 => n9603, B2 => n14613, C1 => n13884, C2 => 
                           n14610, A => n12776, ZN => n12774);
   U11897 : AOI22_X1 port map( A1 => n14607, A2 => n13972, B1 => n14602, B2 => 
                           n14378, ZN => n12776);
   U11898 : OAI221_X1 port map( B1 => n9602, B2 => n14613, C1 => n13885, C2 => 
                           n14610, A => n12759, ZN => n12757);
   U11899 : AOI22_X1 port map( A1 => n14607, A2 => n13973, B1 => n14602, B2 => 
                           n14379, ZN => n12759);
   U11900 : OAI221_X1 port map( B1 => n9601, B2 => n14613, C1 => n13886, C2 => 
                           n14610, A => n12742, ZN => n12740);
   U11901 : AOI22_X1 port map( A1 => n14607, A2 => n13974, B1 => n14602, B2 => 
                           n14380, ZN => n12742);
   U11902 : OAI221_X1 port map( B1 => n9600, B2 => n14613, C1 => n13887, C2 => 
                           n14610, A => n12725, ZN => n12723);
   U11903 : AOI22_X1 port map( A1 => n14607, A2 => n13975, B1 => n14602, B2 => 
                           n14381, ZN => n12725);
   U11904 : OAI221_X1 port map( B1 => n9599, B2 => n14613, C1 => n13888, C2 => 
                           n14610, A => n12708, ZN => n12706);
   U11905 : AOI22_X1 port map( A1 => n14607, A2 => n13976, B1 => n14602, B2 => 
                           n14382, ZN => n12708);
   U11906 : OAI221_X1 port map( B1 => n9598, B2 => n14613, C1 => n13889, C2 => 
                           n14610, A => n12691, ZN => n12689);
   U11907 : AOI22_X1 port map( A1 => n14607, A2 => n13977, B1 => n14602, B2 => 
                           n14383, ZN => n12691);
   U11908 : OAI221_X1 port map( B1 => n9597, B2 => n14613, C1 => n13890, C2 => 
                           n14610, A => n12674, ZN => n12672);
   U11909 : AOI22_X1 port map( A1 => n14607, A2 => n13978, B1 => n14602, B2 => 
                           n14384, ZN => n12674);
   U11910 : OAI221_X1 port map( B1 => n9596, B2 => n14613, C1 => n13891, C2 => 
                           n14610, A => n12649, ZN => n12643);
   U11911 : AOI22_X1 port map( A1 => n14607, A2 => n13979, B1 => n14602, B2 => 
                           n14385, ZN => n12649);
   U11912 : OAI221_X1 port map( B1 => n9603, B2 => n14711, C1 => n13884, C2 => 
                           n14708, A => n12195, ZN => n12193);
   U11913 : AOI22_X1 port map( A1 => n14705, A2 => n13972, B1 => n14700, B2 => 
                           n14378, ZN => n12195);
   U11914 : OAI221_X1 port map( B1 => n9602, B2 => n14711, C1 => n13885, C2 => 
                           n14708, A => n12178, ZN => n12176);
   U11915 : AOI22_X1 port map( A1 => n14705, A2 => n13973, B1 => n14700, B2 => 
                           n14379, ZN => n12178);
   U11916 : OAI221_X1 port map( B1 => n9601, B2 => n14711, C1 => n13886, C2 => 
                           n14708, A => n12161, ZN => n12159);
   U11917 : AOI22_X1 port map( A1 => n14705, A2 => n13974, B1 => n14700, B2 => 
                           n14380, ZN => n12161);
   U11918 : OAI221_X1 port map( B1 => n9600, B2 => n14711, C1 => n13887, C2 => 
                           n14708, A => n12144, ZN => n12142);
   U11919 : AOI22_X1 port map( A1 => n14705, A2 => n13975, B1 => n14700, B2 => 
                           n14381, ZN => n12144);
   U11920 : OAI221_X1 port map( B1 => n9599, B2 => n14711, C1 => n13888, C2 => 
                           n14708, A => n12127, ZN => n12125);
   U11921 : AOI22_X1 port map( A1 => n14705, A2 => n13976, B1 => n14700, B2 => 
                           n14382, ZN => n12127);
   U11922 : OAI221_X1 port map( B1 => n9598, B2 => n14711, C1 => n13889, C2 => 
                           n14708, A => n12110, ZN => n12108);
   U11923 : AOI22_X1 port map( A1 => n14705, A2 => n13977, B1 => n14700, B2 => 
                           n14383, ZN => n12110);
   U11924 : OAI221_X1 port map( B1 => n9597, B2 => n14711, C1 => n13890, C2 => 
                           n14708, A => n12093, ZN => n12091);
   U11925 : AOI22_X1 port map( A1 => n14705, A2 => n13978, B1 => n14700, B2 => 
                           n14384, ZN => n12093);
   U11926 : OAI221_X1 port map( B1 => n9596, B2 => n14711, C1 => n13891, C2 => 
                           n14708, A => n12068, ZN => n12062);
   U11927 : AOI22_X1 port map( A1 => n14705, A2 => n13979, B1 => n14700, B2 => 
                           n14385, ZN => n12068);
   U11928 : OAI22_X1 port map( A1 => n14936, A2 => n15062, B1 => n14935, B2 => 
                           n14530, ZN => n1886);
   U11929 : OAI22_X1 port map( A1 => n14936, A2 => n15065, B1 => n14935, B2 => 
                           n14531, ZN => n1887);
   U11930 : OAI22_X1 port map( A1 => n14936, A2 => n15068, B1 => n14935, B2 => 
                           n14532, ZN => n1888);
   U11931 : OAI22_X1 port map( A1 => n14936, A2 => n15071, B1 => n14935, B2 => 
                           n14533, ZN => n1889);
   U11932 : OAI22_X1 port map( A1 => n14936, A2 => n15074, B1 => n14935, B2 => 
                           n14534, ZN => n1890);
   U11933 : OAI22_X1 port map( A1 => n14937, A2 => n15077, B1 => n14935, B2 => 
                           n14535, ZN => n1891);
   U11934 : OAI22_X1 port map( A1 => n14937, A2 => n15080, B1 => n14935, B2 => 
                           n14536, ZN => n1892);
   U11935 : OAI22_X1 port map( A1 => n14937, A2 => n15083, B1 => n14935, B2 => 
                           n14537, ZN => n1893);
   U11936 : OAI22_X1 port map( A1 => n14937, A2 => n15086, B1 => n14935, B2 => 
                           n14538, ZN => n1894);
   U11937 : OAI22_X1 port map( A1 => n14937, A2 => n15089, B1 => n14935, B2 => 
                           n14539, ZN => n1895);
   U11938 : OAI22_X1 port map( A1 => n14938, A2 => n15092, B1 => n14935, B2 => 
                           n14540, ZN => n1896);
   U11939 : OAI22_X1 port map( A1 => n14938, A2 => n15095, B1 => n14935, B2 => 
                           n14541, ZN => n1897);
   U11940 : OAI22_X1 port map( A1 => n14938, A2 => n15098, B1 => n12003, B2 => 
                           n14542, ZN => n1898);
   U11941 : OAI22_X1 port map( A1 => n14938, A2 => n15101, B1 => n12003, B2 => 
                           n14543, ZN => n1899);
   U11942 : OAI22_X1 port map( A1 => n14938, A2 => n15104, B1 => n12003, B2 => 
                           n14544, ZN => n1900);
   U11943 : OAI22_X1 port map( A1 => n14939, A2 => n15107, B1 => n14935, B2 => 
                           n14545, ZN => n1901);
   U11944 : OAI22_X1 port map( A1 => n14939, A2 => n15110, B1 => n14935, B2 => 
                           n14546, ZN => n1902);
   U11945 : OAI22_X1 port map( A1 => n14939, A2 => n15113, B1 => n14935, B2 => 
                           n14547, ZN => n1903);
   U11946 : OAI22_X1 port map( A1 => n14939, A2 => n15116, B1 => n14935, B2 => 
                           n14548, ZN => n1904);
   U11947 : OAI22_X1 port map( A1 => n14939, A2 => n15119, B1 => n14935, B2 => 
                           n14549, ZN => n1905);
   U11948 : OAI22_X1 port map( A1 => n14940, A2 => n15122, B1 => n14935, B2 => 
                           n14550, ZN => n1906);
   U11949 : OAI22_X1 port map( A1 => n14940, A2 => n15125, B1 => n14935, B2 => 
                           n14551, ZN => n1907);
   U11950 : OAI22_X1 port map( A1 => n14940, A2 => n15128, B1 => n14935, B2 => 
                           n14552, ZN => n1908);
   U11951 : OAI22_X1 port map( A1 => n14940, A2 => n15131, B1 => n14935, B2 => 
                           n14553, ZN => n1909);
   U11952 : OAI22_X1 port map( A1 => n14945, A2 => n15062, B1 => n14944, B2 => 
                           n14410, ZN => n1918);
   U11953 : OAI22_X1 port map( A1 => n14945, A2 => n15065, B1 => n14944, B2 => 
                           n14411, ZN => n1919);
   U11954 : OAI22_X1 port map( A1 => n14945, A2 => n15068, B1 => n14944, B2 => 
                           n14412, ZN => n1920);
   U11955 : OAI22_X1 port map( A1 => n14945, A2 => n15071, B1 => n14944, B2 => 
                           n14413, ZN => n1921);
   U11956 : OAI22_X1 port map( A1 => n14945, A2 => n15074, B1 => n14944, B2 => 
                           n14414, ZN => n1922);
   U11957 : OAI22_X1 port map( A1 => n14946, A2 => n15077, B1 => n14944, B2 => 
                           n14415, ZN => n1923);
   U11958 : OAI22_X1 port map( A1 => n14946, A2 => n15080, B1 => n14944, B2 => 
                           n14416, ZN => n1924);
   U11959 : OAI22_X1 port map( A1 => n14946, A2 => n15083, B1 => n14944, B2 => 
                           n14417, ZN => n1925);
   U11960 : OAI22_X1 port map( A1 => n14946, A2 => n15086, B1 => n14944, B2 => 
                           n14418, ZN => n1926);
   U11961 : OAI22_X1 port map( A1 => n14946, A2 => n15089, B1 => n14944, B2 => 
                           n14419, ZN => n1927);
   U11962 : OAI22_X1 port map( A1 => n14947, A2 => n15092, B1 => n14944, B2 => 
                           n14420, ZN => n1928);
   U11963 : OAI22_X1 port map( A1 => n14947, A2 => n15095, B1 => n14944, B2 => 
                           n14421, ZN => n1929);
   U11964 : OAI22_X1 port map( A1 => n14947, A2 => n15098, B1 => n12002, B2 => 
                           n14422, ZN => n1930);
   U11965 : OAI22_X1 port map( A1 => n14947, A2 => n15101, B1 => n12002, B2 => 
                           n14423, ZN => n1931);
   U11966 : OAI22_X1 port map( A1 => n14947, A2 => n15104, B1 => n12002, B2 => 
                           n14424, ZN => n1932);
   U11967 : OAI22_X1 port map( A1 => n14948, A2 => n15107, B1 => n14944, B2 => 
                           n14425, ZN => n1933);
   U11968 : OAI22_X1 port map( A1 => n14948, A2 => n15110, B1 => n14944, B2 => 
                           n14426, ZN => n1934);
   U11969 : OAI22_X1 port map( A1 => n14948, A2 => n15113, B1 => n14944, B2 => 
                           n14427, ZN => n1935);
   U11970 : OAI22_X1 port map( A1 => n14948, A2 => n15116, B1 => n14944, B2 => 
                           n14428, ZN => n1936);
   U11971 : OAI22_X1 port map( A1 => n14948, A2 => n15119, B1 => n14944, B2 => 
                           n14429, ZN => n1937);
   U11972 : OAI22_X1 port map( A1 => n14949, A2 => n15122, B1 => n14944, B2 => 
                           n14430, ZN => n1938);
   U11973 : OAI22_X1 port map( A1 => n14949, A2 => n15125, B1 => n14944, B2 => 
                           n14431, ZN => n1939);
   U11974 : OAI22_X1 port map( A1 => n14949, A2 => n15128, B1 => n14944, B2 => 
                           n14432, ZN => n1940);
   U11975 : OAI22_X1 port map( A1 => n14949, A2 => n15131, B1 => n14944, B2 => 
                           n14433, ZN => n1941);
   U11976 : OAI22_X1 port map( A1 => n14999, A2 => n15061, B1 => n14998, B2 => 
                           n14434, ZN => n2110);
   U11977 : OAI22_X1 port map( A1 => n14999, A2 => n15064, B1 => n14998, B2 => 
                           n14435, ZN => n2111);
   U11978 : OAI22_X1 port map( A1 => n14999, A2 => n15067, B1 => n14998, B2 => 
                           n14436, ZN => n2112);
   U11979 : OAI22_X1 port map( A1 => n14999, A2 => n15070, B1 => n14998, B2 => 
                           n14437, ZN => n2113);
   U11980 : OAI22_X1 port map( A1 => n14999, A2 => n15073, B1 => n14998, B2 => 
                           n14438, ZN => n2114);
   U11981 : OAI22_X1 port map( A1 => n15000, A2 => n15076, B1 => n14998, B2 => 
                           n14439, ZN => n2115);
   U11982 : OAI22_X1 port map( A1 => n15000, A2 => n15079, B1 => n14998, B2 => 
                           n14440, ZN => n2116);
   U11983 : OAI22_X1 port map( A1 => n15000, A2 => n15082, B1 => n14998, B2 => 
                           n14441, ZN => n2117);
   U11984 : OAI22_X1 port map( A1 => n15000, A2 => n15085, B1 => n14998, B2 => 
                           n14442, ZN => n2118);
   U11985 : OAI22_X1 port map( A1 => n15000, A2 => n15088, B1 => n14998, B2 => 
                           n14443, ZN => n2119);
   U11986 : OAI22_X1 port map( A1 => n15001, A2 => n15091, B1 => n14998, B2 => 
                           n14444, ZN => n2120);
   U11987 : OAI22_X1 port map( A1 => n15001, A2 => n15094, B1 => n14998, B2 => 
                           n14445, ZN => n2121);
   U11988 : OAI22_X1 port map( A1 => n15001, A2 => n15097, B1 => n11994, B2 => 
                           n14446, ZN => n2122);
   U11989 : OAI22_X1 port map( A1 => n15001, A2 => n15100, B1 => n11994, B2 => 
                           n14447, ZN => n2123);
   U11990 : OAI22_X1 port map( A1 => n15001, A2 => n15103, B1 => n11994, B2 => 
                           n14448, ZN => n2124);
   U11991 : OAI22_X1 port map( A1 => n15002, A2 => n15106, B1 => n14998, B2 => 
                           n14449, ZN => n2125);
   U11992 : OAI22_X1 port map( A1 => n15002, A2 => n15109, B1 => n14998, B2 => 
                           n14450, ZN => n2126);
   U11993 : OAI22_X1 port map( A1 => n15002, A2 => n15112, B1 => n14998, B2 => 
                           n14451, ZN => n2127);
   U11994 : OAI22_X1 port map( A1 => n15002, A2 => n15115, B1 => n14998, B2 => 
                           n14452, ZN => n2128);
   U11995 : OAI22_X1 port map( A1 => n15002, A2 => n15118, B1 => n14998, B2 => 
                           n14453, ZN => n2129);
   U11996 : OAI22_X1 port map( A1 => n15003, A2 => n15121, B1 => n14998, B2 => 
                           n14454, ZN => n2130);
   U11997 : OAI22_X1 port map( A1 => n15003, A2 => n15124, B1 => n14998, B2 => 
                           n14455, ZN => n2131);
   U11998 : OAI22_X1 port map( A1 => n15003, A2 => n15127, B1 => n14998, B2 => 
                           n14456, ZN => n2132);
   U11999 : OAI22_X1 port map( A1 => n15003, A2 => n15130, B1 => n14998, B2 => 
                           n14457, ZN => n2133);
   U12000 : OAI22_X1 port map( A1 => n15008, A2 => n15061, B1 => n15007, B2 => 
                           n14554, ZN => n2142);
   U12001 : OAI22_X1 port map( A1 => n15008, A2 => n15064, B1 => n15007, B2 => 
                           n14555, ZN => n2143);
   U12002 : OAI22_X1 port map( A1 => n15008, A2 => n15067, B1 => n15007, B2 => 
                           n14556, ZN => n2144);
   U12003 : OAI22_X1 port map( A1 => n15008, A2 => n15070, B1 => n15007, B2 => 
                           n14557, ZN => n2145);
   U12004 : OAI22_X1 port map( A1 => n15008, A2 => n15073, B1 => n15007, B2 => 
                           n14558, ZN => n2146);
   U12005 : OAI22_X1 port map( A1 => n15009, A2 => n15076, B1 => n15007, B2 => 
                           n14559, ZN => n2147);
   U12006 : OAI22_X1 port map( A1 => n15009, A2 => n15079, B1 => n15007, B2 => 
                           n14560, ZN => n2148);
   U12007 : OAI22_X1 port map( A1 => n15009, A2 => n15082, B1 => n15007, B2 => 
                           n14561, ZN => n2149);
   U12008 : OAI22_X1 port map( A1 => n15009, A2 => n15085, B1 => n15007, B2 => 
                           n14562, ZN => n2150);
   U12009 : OAI22_X1 port map( A1 => n15009, A2 => n15088, B1 => n15007, B2 => 
                           n14563, ZN => n2151);
   U12010 : OAI22_X1 port map( A1 => n15010, A2 => n15091, B1 => n15007, B2 => 
                           n14564, ZN => n2152);
   U12011 : OAI22_X1 port map( A1 => n15010, A2 => n15094, B1 => n15007, B2 => 
                           n14565, ZN => n2153);
   U12012 : OAI22_X1 port map( A1 => n15010, A2 => n15097, B1 => n11993, B2 => 
                           n14566, ZN => n2154);
   U12013 : OAI22_X1 port map( A1 => n15010, A2 => n15100, B1 => n11993, B2 => 
                           n14567, ZN => n2155);
   U12014 : OAI22_X1 port map( A1 => n15010, A2 => n15103, B1 => n11993, B2 => 
                           n14568, ZN => n2156);
   U12015 : OAI22_X1 port map( A1 => n15011, A2 => n15106, B1 => n15007, B2 => 
                           n14569, ZN => n2157);
   U12016 : OAI22_X1 port map( A1 => n15011, A2 => n15109, B1 => n15007, B2 => 
                           n14570, ZN => n2158);
   U12017 : OAI22_X1 port map( A1 => n15011, A2 => n15112, B1 => n15007, B2 => 
                           n14571, ZN => n2159);
   U12018 : OAI22_X1 port map( A1 => n15011, A2 => n15115, B1 => n15007, B2 => 
                           n14572, ZN => n2160);
   U12019 : OAI22_X1 port map( A1 => n15011, A2 => n15118, B1 => n15007, B2 => 
                           n14573, ZN => n2161);
   U12020 : OAI22_X1 port map( A1 => n15012, A2 => n15121, B1 => n15007, B2 => 
                           n14574, ZN => n2162);
   U12021 : OAI22_X1 port map( A1 => n15012, A2 => n15124, B1 => n15007, B2 => 
                           n14575, ZN => n2163);
   U12022 : OAI22_X1 port map( A1 => n15012, A2 => n15127, B1 => n15007, B2 => 
                           n14576, ZN => n2164);
   U12023 : OAI22_X1 port map( A1 => n15012, A2 => n15130, B1 => n15007, B2 => 
                           n14577, ZN => n2165);
   U12024 : OAI22_X1 port map( A1 => n15017, A2 => n15061, B1 => n15016, B2 => 
                           n14386, ZN => n2174);
   U12025 : OAI22_X1 port map( A1 => n15017, A2 => n15064, B1 => n15016, B2 => 
                           n14387, ZN => n2175);
   U12026 : OAI22_X1 port map( A1 => n15017, A2 => n15067, B1 => n15016, B2 => 
                           n14388, ZN => n2176);
   U12027 : OAI22_X1 port map( A1 => n15017, A2 => n15070, B1 => n15016, B2 => 
                           n14389, ZN => n2177);
   U12028 : OAI22_X1 port map( A1 => n15017, A2 => n15073, B1 => n15016, B2 => 
                           n14390, ZN => n2178);
   U12029 : OAI22_X1 port map( A1 => n15018, A2 => n15076, B1 => n15016, B2 => 
                           n14391, ZN => n2179);
   U12030 : OAI22_X1 port map( A1 => n15018, A2 => n15079, B1 => n15016, B2 => 
                           n14392, ZN => n2180);
   U12031 : OAI22_X1 port map( A1 => n15018, A2 => n15082, B1 => n15016, B2 => 
                           n14393, ZN => n2181);
   U12032 : OAI22_X1 port map( A1 => n15018, A2 => n15085, B1 => n15016, B2 => 
                           n14394, ZN => n2182);
   U12033 : OAI22_X1 port map( A1 => n15018, A2 => n15088, B1 => n15016, B2 => 
                           n14395, ZN => n2183);
   U12034 : OAI22_X1 port map( A1 => n15019, A2 => n15091, B1 => n15016, B2 => 
                           n14396, ZN => n2184);
   U12035 : OAI22_X1 port map( A1 => n15019, A2 => n15094, B1 => n15016, B2 => 
                           n14397, ZN => n2185);
   U12036 : OAI22_X1 port map( A1 => n15019, A2 => n15097, B1 => n11992, B2 => 
                           n14398, ZN => n2186);
   U12037 : OAI22_X1 port map( A1 => n15019, A2 => n15100, B1 => n11992, B2 => 
                           n14399, ZN => n2187);
   U12038 : OAI22_X1 port map( A1 => n15019, A2 => n15103, B1 => n11992, B2 => 
                           n14400, ZN => n2188);
   U12039 : OAI22_X1 port map( A1 => n15020, A2 => n15106, B1 => n15016, B2 => 
                           n14401, ZN => n2189);
   U12040 : OAI22_X1 port map( A1 => n15020, A2 => n15109, B1 => n15016, B2 => 
                           n14402, ZN => n2190);
   U12041 : OAI22_X1 port map( A1 => n15020, A2 => n15112, B1 => n15016, B2 => 
                           n14403, ZN => n2191);
   U12042 : OAI22_X1 port map( A1 => n15020, A2 => n15115, B1 => n15016, B2 => 
                           n14404, ZN => n2192);
   U12043 : OAI22_X1 port map( A1 => n15020, A2 => n15118, B1 => n15016, B2 => 
                           n14405, ZN => n2193);
   U12044 : OAI22_X1 port map( A1 => n15021, A2 => n15121, B1 => n15016, B2 => 
                           n14406, ZN => n2194);
   U12045 : OAI22_X1 port map( A1 => n15021, A2 => n15124, B1 => n15016, B2 => 
                           n14407, ZN => n2195);
   U12046 : OAI22_X1 port map( A1 => n15021, A2 => n15127, B1 => n15016, B2 => 
                           n14408, ZN => n2196);
   U12047 : OAI22_X1 port map( A1 => n15021, A2 => n15130, B1 => n15016, B2 => 
                           n14409, ZN => n2197);
   U12048 : OAI22_X1 port map( A1 => n15035, A2 => n15061, B1 => n15034, B2 => 
                           n14458, ZN => n2238);
   U12049 : OAI22_X1 port map( A1 => n15035, A2 => n15064, B1 => n15034, B2 => 
                           n14459, ZN => n2239);
   U12050 : OAI22_X1 port map( A1 => n15035, A2 => n15067, B1 => n15034, B2 => 
                           n14460, ZN => n2240);
   U12051 : OAI22_X1 port map( A1 => n15035, A2 => n15070, B1 => n15034, B2 => 
                           n14461, ZN => n2241);
   U12052 : OAI22_X1 port map( A1 => n15035, A2 => n15073, B1 => n15034, B2 => 
                           n14462, ZN => n2242);
   U12053 : OAI22_X1 port map( A1 => n15036, A2 => n15076, B1 => n15034, B2 => 
                           n14463, ZN => n2243);
   U12054 : OAI22_X1 port map( A1 => n15036, A2 => n15079, B1 => n15034, B2 => 
                           n14464, ZN => n2244);
   U12055 : OAI22_X1 port map( A1 => n15036, A2 => n15082, B1 => n15034, B2 => 
                           n14465, ZN => n2245);
   U12056 : OAI22_X1 port map( A1 => n15036, A2 => n15085, B1 => n15034, B2 => 
                           n14466, ZN => n2246);
   U12057 : OAI22_X1 port map( A1 => n15036, A2 => n15088, B1 => n15034, B2 => 
                           n14467, ZN => n2247);
   U12058 : OAI22_X1 port map( A1 => n15037, A2 => n15091, B1 => n15034, B2 => 
                           n14468, ZN => n2248);
   U12059 : OAI22_X1 port map( A1 => n15037, A2 => n15094, B1 => n15034, B2 => 
                           n14469, ZN => n2249);
   U12060 : OAI22_X1 port map( A1 => n15037, A2 => n15097, B1 => n11987, B2 => 
                           n14470, ZN => n2250);
   U12061 : OAI22_X1 port map( A1 => n15037, A2 => n15100, B1 => n11987, B2 => 
                           n14471, ZN => n2251);
   U12062 : OAI22_X1 port map( A1 => n15037, A2 => n15103, B1 => n11987, B2 => 
                           n14472, ZN => n2252);
   U12063 : OAI22_X1 port map( A1 => n15038, A2 => n15106, B1 => n15034, B2 => 
                           n14473, ZN => n2253);
   U12064 : OAI22_X1 port map( A1 => n15038, A2 => n15109, B1 => n15034, B2 => 
                           n14474, ZN => n2254);
   U12065 : OAI22_X1 port map( A1 => n15038, A2 => n15112, B1 => n15034, B2 => 
                           n14475, ZN => n2255);
   U12066 : OAI22_X1 port map( A1 => n15038, A2 => n15115, B1 => n15034, B2 => 
                           n14476, ZN => n2256);
   U12067 : OAI22_X1 port map( A1 => n15038, A2 => n15118, B1 => n15034, B2 => 
                           n14477, ZN => n2257);
   U12068 : OAI22_X1 port map( A1 => n15039, A2 => n15121, B1 => n15034, B2 => 
                           n14478, ZN => n2258);
   U12069 : OAI22_X1 port map( A1 => n15039, A2 => n15124, B1 => n15034, B2 => 
                           n14479, ZN => n2259);
   U12070 : OAI22_X1 port map( A1 => n15039, A2 => n15127, B1 => n15034, B2 => 
                           n14480, ZN => n2260);
   U12071 : OAI22_X1 port map( A1 => n15039, A2 => n15130, B1 => n15034, B2 => 
                           n14481, ZN => n2261);
   U12072 : OAI22_X1 port map( A1 => n9659, A2 => n12025, B1 => n14781, B2 => 
                           n15063, ZN => n1342);
   U12073 : OAI22_X1 port map( A1 => n9648, A2 => n14780, B1 => n14783, B2 => 
                           n15096, ZN => n1353);
   U12074 : OAI22_X1 port map( A1 => n9647, A2 => n14780, B1 => n14784, B2 => 
                           n15099, ZN => n1354);
   U12075 : OAI22_X1 port map( A1 => n9646, A2 => n14780, B1 => n14784, B2 => 
                           n15102, ZN => n1355);
   U12076 : OAI22_X1 port map( A1 => n9645, A2 => n14780, B1 => n14784, B2 => 
                           n15105, ZN => n1356);
   U12077 : OAI22_X1 port map( A1 => n9644, A2 => n14780, B1 => n14784, B2 => 
                           n15108, ZN => n1357);
   U12078 : OAI22_X1 port map( A1 => n9643, A2 => n14780, B1 => n14785, B2 => 
                           n15111, ZN => n1358);
   U12079 : OAI22_X1 port map( A1 => n9642, A2 => n14780, B1 => n14785, B2 => 
                           n15114, ZN => n1359);
   U12080 : OAI22_X1 port map( A1 => n9641, A2 => n14780, B1 => n14785, B2 => 
                           n15117, ZN => n1360);
   U12081 : OAI22_X1 port map( A1 => n9640, A2 => n14780, B1 => n14785, B2 => 
                           n15120, ZN => n1361);
   U12082 : OAI22_X1 port map( A1 => n9639, A2 => n12025, B1 => n14786, B2 => 
                           n15123, ZN => n1362);
   U12083 : OAI22_X1 port map( A1 => n9638, A2 => n14780, B1 => n14786, B2 => 
                           n15126, ZN => n1363);
   U12084 : OAI22_X1 port map( A1 => n9637, A2 => n12025, B1 => n14786, B2 => 
                           n15129, ZN => n1364);
   U12085 : OAI22_X1 port map( A1 => n9636, A2 => n14780, B1 => n14786, B2 => 
                           n15132, ZN => n1365);
   U12086 : OAI22_X1 port map( A1 => n9635, A2 => n12025, B1 => n14787, B2 => 
                           n15135, ZN => n1366);
   U12087 : OAI22_X1 port map( A1 => n9634, A2 => n14780, B1 => n14787, B2 => 
                           n15138, ZN => n1367);
   U12088 : OAI22_X1 port map( A1 => n9633, A2 => n12025, B1 => n14787, B2 => 
                           n15141, ZN => n1368);
   U12089 : OAI22_X1 port map( A1 => n9632, A2 => n14780, B1 => n14787, B2 => 
                           n15144, ZN => n1369);
   U12090 : OAI22_X1 port map( A1 => n9631, A2 => n12025, B1 => n14788, B2 => 
                           n15147, ZN => n1370);
   U12091 : OAI22_X1 port map( A1 => n9630, A2 => n14780, B1 => n14788, B2 => 
                           n15150, ZN => n1371);
   U12092 : OAI22_X1 port map( A1 => n14792, A2 => n15063, B1 => n9627, B2 => 
                           n14791, ZN => n1374);
   U12093 : OAI22_X1 port map( A1 => n14792, A2 => n15066, B1 => n9626, B2 => 
                           n14791, ZN => n1375);
   U12094 : OAI22_X1 port map( A1 => n14792, A2 => n15069, B1 => n9625, B2 => 
                           n14791, ZN => n1376);
   U12095 : OAI22_X1 port map( A1 => n14792, A2 => n15072, B1 => n9624, B2 => 
                           n14791, ZN => n1377);
   U12096 : OAI22_X1 port map( A1 => n14792, A2 => n15075, B1 => n9623, B2 => 
                           n14791, ZN => n1378);
   U12097 : OAI22_X1 port map( A1 => n14793, A2 => n15078, B1 => n9622, B2 => 
                           n14791, ZN => n1379);
   U12098 : OAI22_X1 port map( A1 => n14793, A2 => n15081, B1 => n9621, B2 => 
                           n14791, ZN => n1380);
   U12099 : OAI22_X1 port map( A1 => n14793, A2 => n15084, B1 => n9620, B2 => 
                           n14791, ZN => n1381);
   U12100 : OAI22_X1 port map( A1 => n14793, A2 => n15087, B1 => n9619, B2 => 
                           n14791, ZN => n1382);
   U12101 : OAI22_X1 port map( A1 => n14793, A2 => n15090, B1 => n9618, B2 => 
                           n14791, ZN => n1383);
   U12102 : OAI22_X1 port map( A1 => n14794, A2 => n15093, B1 => n9617, B2 => 
                           n14791, ZN => n1384);
   U12103 : OAI22_X1 port map( A1 => n14794, A2 => n15096, B1 => n9616, B2 => 
                           n14791, ZN => n1385);
   U12104 : OAI22_X1 port map( A1 => n14794, A2 => n15099, B1 => n9615, B2 => 
                           n12024, ZN => n1386);
   U12105 : OAI22_X1 port map( A1 => n14794, A2 => n15102, B1 => n9614, B2 => 
                           n12024, ZN => n1387);
   U12106 : OAI22_X1 port map( A1 => n14794, A2 => n15105, B1 => n9613, B2 => 
                           n12024, ZN => n1388);
   U12107 : OAI22_X1 port map( A1 => n14795, A2 => n15108, B1 => n9612, B2 => 
                           n14791, ZN => n1389);
   U12108 : OAI22_X1 port map( A1 => n14795, A2 => n15111, B1 => n9611, B2 => 
                           n14791, ZN => n1390);
   U12109 : OAI22_X1 port map( A1 => n14795, A2 => n15114, B1 => n9610, B2 => 
                           n14791, ZN => n1391);
   U12110 : OAI22_X1 port map( A1 => n14795, A2 => n15117, B1 => n9609, B2 => 
                           n14791, ZN => n1392);
   U12111 : OAI22_X1 port map( A1 => n14795, A2 => n15120, B1 => n9608, B2 => 
                           n14791, ZN => n1393);
   U12112 : OAI22_X1 port map( A1 => n14796, A2 => n15123, B1 => n9607, B2 => 
                           n14791, ZN => n1394);
   U12113 : OAI22_X1 port map( A1 => n14796, A2 => n15126, B1 => n9606, B2 => 
                           n14791, ZN => n1395);
   U12114 : OAI22_X1 port map( A1 => n14796, A2 => n15129, B1 => n9605, B2 => 
                           n14791, ZN => n1396);
   U12115 : OAI22_X1 port map( A1 => n14796, A2 => n15132, B1 => n9604, B2 => 
                           n14791, ZN => n1397);
   U12116 : OAI22_X1 port map( A1 => n14819, A2 => n15063, B1 => n9531, B2 => 
                           n14818, ZN => n1470);
   U12117 : OAI22_X1 port map( A1 => n14819, A2 => n15066, B1 => n9530, B2 => 
                           n14818, ZN => n1471);
   U12118 : OAI22_X1 port map( A1 => n14819, A2 => n15069, B1 => n9529, B2 => 
                           n14818, ZN => n1472);
   U12119 : OAI22_X1 port map( A1 => n14819, A2 => n15072, B1 => n9528, B2 => 
                           n14818, ZN => n1473);
   U12120 : OAI22_X1 port map( A1 => n14819, A2 => n15075, B1 => n9527, B2 => 
                           n14818, ZN => n1474);
   U12121 : OAI22_X1 port map( A1 => n14820, A2 => n15078, B1 => n9526, B2 => 
                           n14818, ZN => n1475);
   U12122 : OAI22_X1 port map( A1 => n14820, A2 => n15081, B1 => n9525, B2 => 
                           n14818, ZN => n1476);
   U12123 : OAI22_X1 port map( A1 => n14820, A2 => n15084, B1 => n9524, B2 => 
                           n14818, ZN => n1477);
   U12124 : OAI22_X1 port map( A1 => n14820, A2 => n15087, B1 => n9523, B2 => 
                           n14818, ZN => n1478);
   U12125 : OAI22_X1 port map( A1 => n14820, A2 => n15090, B1 => n9522, B2 => 
                           n14818, ZN => n1479);
   U12126 : OAI22_X1 port map( A1 => n14821, A2 => n15093, B1 => n9521, B2 => 
                           n14818, ZN => n1480);
   U12127 : OAI22_X1 port map( A1 => n14821, A2 => n15096, B1 => n9520, B2 => 
                           n14818, ZN => n1481);
   U12128 : OAI22_X1 port map( A1 => n14821, A2 => n15099, B1 => n9519, B2 => 
                           n12020, ZN => n1482);
   U12129 : OAI22_X1 port map( A1 => n14821, A2 => n15102, B1 => n9518, B2 => 
                           n12020, ZN => n1483);
   U12130 : OAI22_X1 port map( A1 => n14821, A2 => n15105, B1 => n9517, B2 => 
                           n12020, ZN => n1484);
   U12131 : OAI22_X1 port map( A1 => n14822, A2 => n15108, B1 => n9516, B2 => 
                           n14818, ZN => n1485);
   U12132 : OAI22_X1 port map( A1 => n14822, A2 => n15111, B1 => n9515, B2 => 
                           n14818, ZN => n1486);
   U12133 : OAI22_X1 port map( A1 => n14822, A2 => n15114, B1 => n9514, B2 => 
                           n14818, ZN => n1487);
   U12134 : OAI22_X1 port map( A1 => n14822, A2 => n15117, B1 => n9513, B2 => 
                           n14818, ZN => n1488);
   U12135 : OAI22_X1 port map( A1 => n14822, A2 => n15120, B1 => n9512, B2 => 
                           n14818, ZN => n1489);
   U12136 : OAI22_X1 port map( A1 => n14823, A2 => n15123, B1 => n9511, B2 => 
                           n14818, ZN => n1490);
   U12137 : OAI22_X1 port map( A1 => n14823, A2 => n15126, B1 => n9510, B2 => 
                           n14818, ZN => n1491);
   U12138 : OAI22_X1 port map( A1 => n14823, A2 => n15129, B1 => n9509, B2 => 
                           n14818, ZN => n1492);
   U12139 : OAI22_X1 port map( A1 => n14823, A2 => n15132, B1 => n9508, B2 => 
                           n14818, ZN => n1493);
   U12140 : OAI22_X1 port map( A1 => n14801, A2 => n15063, B1 => n9595, B2 => 
                           n14800, ZN => n1406);
   U12141 : OAI22_X1 port map( A1 => n14801, A2 => n15066, B1 => n9594, B2 => 
                           n14800, ZN => n1407);
   U12142 : OAI22_X1 port map( A1 => n14801, A2 => n15069, B1 => n9593, B2 => 
                           n14800, ZN => n1408);
   U12143 : OAI22_X1 port map( A1 => n14801, A2 => n15072, B1 => n9592, B2 => 
                           n14800, ZN => n1409);
   U12144 : OAI22_X1 port map( A1 => n14801, A2 => n15075, B1 => n9591, B2 => 
                           n14800, ZN => n1410);
   U12145 : OAI22_X1 port map( A1 => n14802, A2 => n15078, B1 => n9590, B2 => 
                           n14800, ZN => n1411);
   U12146 : OAI22_X1 port map( A1 => n14802, A2 => n15081, B1 => n9589, B2 => 
                           n14800, ZN => n1412);
   U12147 : OAI22_X1 port map( A1 => n14802, A2 => n15084, B1 => n9588, B2 => 
                           n14800, ZN => n1413);
   U12148 : OAI22_X1 port map( A1 => n14802, A2 => n15087, B1 => n9587, B2 => 
                           n14800, ZN => n1414);
   U12149 : OAI22_X1 port map( A1 => n14802, A2 => n15090, B1 => n9586, B2 => 
                           n14800, ZN => n1415);
   U12150 : OAI22_X1 port map( A1 => n14803, A2 => n15093, B1 => n9585, B2 => 
                           n14800, ZN => n1416);
   U12151 : OAI22_X1 port map( A1 => n14803, A2 => n15096, B1 => n9584, B2 => 
                           n14800, ZN => n1417);
   U12152 : OAI22_X1 port map( A1 => n14803, A2 => n15099, B1 => n9583, B2 => 
                           n12023, ZN => n1418);
   U12153 : OAI22_X1 port map( A1 => n14803, A2 => n15102, B1 => n9582, B2 => 
                           n12023, ZN => n1419);
   U12154 : OAI22_X1 port map( A1 => n14803, A2 => n15105, B1 => n9581, B2 => 
                           n12023, ZN => n1420);
   U12155 : OAI22_X1 port map( A1 => n14804, A2 => n15108, B1 => n9580, B2 => 
                           n14800, ZN => n1421);
   U12156 : OAI22_X1 port map( A1 => n14804, A2 => n15111, B1 => n9579, B2 => 
                           n14800, ZN => n1422);
   U12157 : OAI22_X1 port map( A1 => n14804, A2 => n15114, B1 => n9578, B2 => 
                           n14800, ZN => n1423);
   U12158 : OAI22_X1 port map( A1 => n14804, A2 => n15117, B1 => n9577, B2 => 
                           n14800, ZN => n1424);
   U12159 : OAI22_X1 port map( A1 => n14804, A2 => n15120, B1 => n9576, B2 => 
                           n14800, ZN => n1425);
   U12160 : OAI22_X1 port map( A1 => n14805, A2 => n15123, B1 => n9575, B2 => 
                           n14800, ZN => n1426);
   U12161 : OAI22_X1 port map( A1 => n14805, A2 => n15126, B1 => n9574, B2 => 
                           n14800, ZN => n1427);
   U12162 : OAI22_X1 port map( A1 => n14805, A2 => n15129, B1 => n9573, B2 => 
                           n14800, ZN => n1428);
   U12163 : OAI22_X1 port map( A1 => n14805, A2 => n15132, B1 => n9572, B2 => 
                           n14800, ZN => n1429);
   U12164 : OAI22_X1 port map( A1 => n14810, A2 => n15063, B1 => n9563, B2 => 
                           n14809, ZN => n1438);
   U12165 : OAI22_X1 port map( A1 => n14810, A2 => n15066, B1 => n9562, B2 => 
                           n14809, ZN => n1439);
   U12166 : OAI22_X1 port map( A1 => n14810, A2 => n15069, B1 => n9561, B2 => 
                           n14809, ZN => n1440);
   U12167 : OAI22_X1 port map( A1 => n14810, A2 => n15072, B1 => n9560, B2 => 
                           n14809, ZN => n1441);
   U12168 : OAI22_X1 port map( A1 => n14810, A2 => n15075, B1 => n9559, B2 => 
                           n14809, ZN => n1442);
   U12169 : OAI22_X1 port map( A1 => n14811, A2 => n15078, B1 => n9558, B2 => 
                           n14809, ZN => n1443);
   U12170 : OAI22_X1 port map( A1 => n14811, A2 => n15081, B1 => n9557, B2 => 
                           n14809, ZN => n1444);
   U12171 : OAI22_X1 port map( A1 => n14811, A2 => n15084, B1 => n9556, B2 => 
                           n14809, ZN => n1445);
   U12172 : OAI22_X1 port map( A1 => n14811, A2 => n15087, B1 => n9555, B2 => 
                           n14809, ZN => n1446);
   U12173 : OAI22_X1 port map( A1 => n14811, A2 => n15090, B1 => n9554, B2 => 
                           n14809, ZN => n1447);
   U12174 : OAI22_X1 port map( A1 => n14812, A2 => n15093, B1 => n9553, B2 => 
                           n14809, ZN => n1448);
   U12175 : OAI22_X1 port map( A1 => n14812, A2 => n15096, B1 => n9552, B2 => 
                           n14809, ZN => n1449);
   U12176 : OAI22_X1 port map( A1 => n14812, A2 => n15099, B1 => n9551, B2 => 
                           n12021, ZN => n1450);
   U12177 : OAI22_X1 port map( A1 => n14812, A2 => n15102, B1 => n9550, B2 => 
                           n12021, ZN => n1451);
   U12178 : OAI22_X1 port map( A1 => n14812, A2 => n15105, B1 => n9549, B2 => 
                           n12021, ZN => n1452);
   U12179 : OAI22_X1 port map( A1 => n14813, A2 => n15108, B1 => n9548, B2 => 
                           n14809, ZN => n1453);
   U12180 : OAI22_X1 port map( A1 => n14813, A2 => n15111, B1 => n9547, B2 => 
                           n14809, ZN => n1454);
   U12181 : OAI22_X1 port map( A1 => n14813, A2 => n15114, B1 => n9546, B2 => 
                           n14809, ZN => n1455);
   U12182 : OAI22_X1 port map( A1 => n14813, A2 => n15117, B1 => n9545, B2 => 
                           n14809, ZN => n1456);
   U12183 : OAI22_X1 port map( A1 => n14813, A2 => n15120, B1 => n9544, B2 => 
                           n14809, ZN => n1457);
   U12184 : OAI22_X1 port map( A1 => n14814, A2 => n15123, B1 => n9543, B2 => 
                           n14809, ZN => n1458);
   U12185 : OAI22_X1 port map( A1 => n14814, A2 => n15126, B1 => n9542, B2 => 
                           n14809, ZN => n1459);
   U12186 : OAI22_X1 port map( A1 => n14814, A2 => n15129, B1 => n9541, B2 => 
                           n14809, ZN => n1460);
   U12187 : OAI22_X1 port map( A1 => n14814, A2 => n15132, B1 => n9540, B2 => 
                           n14809, ZN => n1461);
   U12188 : OAI22_X1 port map( A1 => n14828, A2 => n15063, B1 => n9499, B2 => 
                           n14827, ZN => n1502);
   U12189 : OAI22_X1 port map( A1 => n14828, A2 => n15066, B1 => n9498, B2 => 
                           n14827, ZN => n1503);
   U12190 : OAI22_X1 port map( A1 => n14828, A2 => n15069, B1 => n9497, B2 => 
                           n14827, ZN => n1504);
   U12191 : OAI22_X1 port map( A1 => n14828, A2 => n15072, B1 => n9496, B2 => 
                           n14827, ZN => n1505);
   U12192 : OAI22_X1 port map( A1 => n14828, A2 => n15075, B1 => n9495, B2 => 
                           n14827, ZN => n1506);
   U12193 : OAI22_X1 port map( A1 => n14829, A2 => n15078, B1 => n9494, B2 => 
                           n14827, ZN => n1507);
   U12194 : OAI22_X1 port map( A1 => n14829, A2 => n15081, B1 => n9493, B2 => 
                           n14827, ZN => n1508);
   U12195 : OAI22_X1 port map( A1 => n14829, A2 => n15084, B1 => n9492, B2 => 
                           n14827, ZN => n1509);
   U12196 : OAI22_X1 port map( A1 => n14829, A2 => n15087, B1 => n9491, B2 => 
                           n14827, ZN => n1510);
   U12197 : OAI22_X1 port map( A1 => n14829, A2 => n15090, B1 => n9490, B2 => 
                           n14827, ZN => n1511);
   U12198 : OAI22_X1 port map( A1 => n14830, A2 => n15093, B1 => n9489, B2 => 
                           n14827, ZN => n1512);
   U12199 : OAI22_X1 port map( A1 => n14830, A2 => n15096, B1 => n9488, B2 => 
                           n14827, ZN => n1513);
   U12200 : OAI22_X1 port map( A1 => n14830, A2 => n15099, B1 => n9487, B2 => 
                           n12019, ZN => n1514);
   U12201 : OAI22_X1 port map( A1 => n14830, A2 => n15102, B1 => n9486, B2 => 
                           n12019, ZN => n1515);
   U12202 : OAI22_X1 port map( A1 => n14830, A2 => n15105, B1 => n9485, B2 => 
                           n12019, ZN => n1516);
   U12203 : OAI22_X1 port map( A1 => n14831, A2 => n15108, B1 => n9484, B2 => 
                           n14827, ZN => n1517);
   U12204 : OAI22_X1 port map( A1 => n14831, A2 => n15111, B1 => n9483, B2 => 
                           n14827, ZN => n1518);
   U12205 : OAI22_X1 port map( A1 => n14831, A2 => n15114, B1 => n9482, B2 => 
                           n14827, ZN => n1519);
   U12206 : OAI22_X1 port map( A1 => n14831, A2 => n15117, B1 => n9481, B2 => 
                           n14827, ZN => n1520);
   U12207 : OAI22_X1 port map( A1 => n14831, A2 => n15120, B1 => n9480, B2 => 
                           n14827, ZN => n1521);
   U12208 : OAI22_X1 port map( A1 => n14832, A2 => n15123, B1 => n9479, B2 => 
                           n14827, ZN => n1522);
   U12209 : OAI22_X1 port map( A1 => n14832, A2 => n15126, B1 => n9478, B2 => 
                           n14827, ZN => n1523);
   U12210 : OAI22_X1 port map( A1 => n14832, A2 => n15129, B1 => n9477, B2 => 
                           n14827, ZN => n1524);
   U12211 : OAI22_X1 port map( A1 => n14832, A2 => n15132, B1 => n9476, B2 => 
                           n14827, ZN => n1525);
   U12212 : OAI22_X1 port map( A1 => n14837, A2 => n15063, B1 => n9467, B2 => 
                           n14836, ZN => n1534);
   U12213 : OAI22_X1 port map( A1 => n14837, A2 => n15066, B1 => n9466, B2 => 
                           n14836, ZN => n1535);
   U12214 : OAI22_X1 port map( A1 => n14837, A2 => n15069, B1 => n9465, B2 => 
                           n14836, ZN => n1536);
   U12215 : OAI22_X1 port map( A1 => n14837, A2 => n15072, B1 => n9464, B2 => 
                           n14836, ZN => n1537);
   U12216 : OAI22_X1 port map( A1 => n14837, A2 => n15075, B1 => n9463, B2 => 
                           n14836, ZN => n1538);
   U12217 : OAI22_X1 port map( A1 => n14838, A2 => n15078, B1 => n9462, B2 => 
                           n14836, ZN => n1539);
   U12218 : OAI22_X1 port map( A1 => n14838, A2 => n15081, B1 => n9461, B2 => 
                           n14836, ZN => n1540);
   U12219 : OAI22_X1 port map( A1 => n14838, A2 => n15084, B1 => n9460, B2 => 
                           n14836, ZN => n1541);
   U12220 : OAI22_X1 port map( A1 => n14838, A2 => n15087, B1 => n9459, B2 => 
                           n14836, ZN => n1542);
   U12221 : OAI22_X1 port map( A1 => n14838, A2 => n15090, B1 => n9458, B2 => 
                           n14836, ZN => n1543);
   U12222 : OAI22_X1 port map( A1 => n14839, A2 => n15093, B1 => n9457, B2 => 
                           n14836, ZN => n1544);
   U12223 : OAI22_X1 port map( A1 => n14839, A2 => n15096, B1 => n9456, B2 => 
                           n14836, ZN => n1545);
   U12224 : OAI22_X1 port map( A1 => n14839, A2 => n15099, B1 => n9455, B2 => 
                           n12018, ZN => n1546);
   U12225 : OAI22_X1 port map( A1 => n14839, A2 => n15102, B1 => n9454, B2 => 
                           n12018, ZN => n1547);
   U12226 : OAI22_X1 port map( A1 => n14839, A2 => n15105, B1 => n9453, B2 => 
                           n12018, ZN => n1548);
   U12227 : OAI22_X1 port map( A1 => n14840, A2 => n15108, B1 => n9452, B2 => 
                           n14836, ZN => n1549);
   U12228 : OAI22_X1 port map( A1 => n14840, A2 => n15111, B1 => n9451, B2 => 
                           n14836, ZN => n1550);
   U12229 : OAI22_X1 port map( A1 => n14840, A2 => n15114, B1 => n9450, B2 => 
                           n14836, ZN => n1551);
   U12230 : OAI22_X1 port map( A1 => n14840, A2 => n15117, B1 => n9449, B2 => 
                           n14836, ZN => n1552);
   U12231 : OAI22_X1 port map( A1 => n14840, A2 => n15120, B1 => n9448, B2 => 
                           n14836, ZN => n1553);
   U12232 : OAI22_X1 port map( A1 => n14841, A2 => n15123, B1 => n9447, B2 => 
                           n14836, ZN => n1554);
   U12233 : OAI22_X1 port map( A1 => n14841, A2 => n15126, B1 => n9446, B2 => 
                           n14836, ZN => n1555);
   U12234 : OAI22_X1 port map( A1 => n14841, A2 => n15129, B1 => n9445, B2 => 
                           n14836, ZN => n1556);
   U12235 : OAI22_X1 port map( A1 => n14841, A2 => n15132, B1 => n9444, B2 => 
                           n14836, ZN => n1557);
   U12236 : OAI22_X1 port map( A1 => n14846, A2 => n15063, B1 => n9435, B2 => 
                           n14845, ZN => n1566);
   U12237 : OAI22_X1 port map( A1 => n14846, A2 => n15066, B1 => n9434, B2 => 
                           n14845, ZN => n1567);
   U12238 : OAI22_X1 port map( A1 => n14846, A2 => n15069, B1 => n9433, B2 => 
                           n14845, ZN => n1568);
   U12239 : OAI22_X1 port map( A1 => n14846, A2 => n15072, B1 => n9432, B2 => 
                           n14845, ZN => n1569);
   U12240 : OAI22_X1 port map( A1 => n14846, A2 => n15075, B1 => n9431, B2 => 
                           n14845, ZN => n1570);
   U12241 : OAI22_X1 port map( A1 => n14847, A2 => n15078, B1 => n9430, B2 => 
                           n14845, ZN => n1571);
   U12242 : OAI22_X1 port map( A1 => n14847, A2 => n15081, B1 => n9429, B2 => 
                           n14845, ZN => n1572);
   U12243 : OAI22_X1 port map( A1 => n14847, A2 => n15084, B1 => n9428, B2 => 
                           n14845, ZN => n1573);
   U12244 : OAI22_X1 port map( A1 => n14847, A2 => n15087, B1 => n9427, B2 => 
                           n14845, ZN => n1574);
   U12245 : OAI22_X1 port map( A1 => n14847, A2 => n15090, B1 => n9426, B2 => 
                           n14845, ZN => n1575);
   U12246 : OAI22_X1 port map( A1 => n14848, A2 => n15093, B1 => n9425, B2 => 
                           n14845, ZN => n1576);
   U12247 : OAI22_X1 port map( A1 => n14848, A2 => n15096, B1 => n9424, B2 => 
                           n14845, ZN => n1577);
   U12248 : OAI22_X1 port map( A1 => n14848, A2 => n15099, B1 => n9423, B2 => 
                           n12016, ZN => n1578);
   U12249 : OAI22_X1 port map( A1 => n14848, A2 => n15102, B1 => n9422, B2 => 
                           n12016, ZN => n1579);
   U12250 : OAI22_X1 port map( A1 => n14848, A2 => n15105, B1 => n9421, B2 => 
                           n12016, ZN => n1580);
   U12251 : OAI22_X1 port map( A1 => n14849, A2 => n15108, B1 => n9420, B2 => 
                           n14845, ZN => n1581);
   U12252 : OAI22_X1 port map( A1 => n14849, A2 => n15111, B1 => n9419, B2 => 
                           n14845, ZN => n1582);
   U12253 : OAI22_X1 port map( A1 => n14849, A2 => n15114, B1 => n9418, B2 => 
                           n14845, ZN => n1583);
   U12254 : OAI22_X1 port map( A1 => n14849, A2 => n15117, B1 => n9417, B2 => 
                           n14845, ZN => n1584);
   U12255 : OAI22_X1 port map( A1 => n14849, A2 => n15120, B1 => n9416, B2 => 
                           n14845, ZN => n1585);
   U12256 : OAI22_X1 port map( A1 => n14850, A2 => n15123, B1 => n9415, B2 => 
                           n14845, ZN => n1586);
   U12257 : OAI22_X1 port map( A1 => n14850, A2 => n15126, B1 => n9414, B2 => 
                           n14845, ZN => n1587);
   U12258 : OAI22_X1 port map( A1 => n14850, A2 => n15129, B1 => n9413, B2 => 
                           n14845, ZN => n1588);
   U12259 : OAI22_X1 port map( A1 => n14850, A2 => n15132, B1 => n9412, B2 => 
                           n14845, ZN => n1589);
   U12260 : OAI22_X1 port map( A1 => n14927, A2 => n15062, B1 => n9147, B2 => 
                           n14926, ZN => n1854);
   U12261 : OAI22_X1 port map( A1 => n14927, A2 => n15065, B1 => n9146, B2 => 
                           n14926, ZN => n1855);
   U12262 : OAI22_X1 port map( A1 => n14927, A2 => n15068, B1 => n9145, B2 => 
                           n14926, ZN => n1856);
   U12263 : OAI22_X1 port map( A1 => n14927, A2 => n15071, B1 => n9144, B2 => 
                           n14926, ZN => n1857);
   U12264 : OAI22_X1 port map( A1 => n14927, A2 => n15074, B1 => n9143, B2 => 
                           n14926, ZN => n1858);
   U12265 : OAI22_X1 port map( A1 => n14928, A2 => n15077, B1 => n9142, B2 => 
                           n14926, ZN => n1859);
   U12266 : OAI22_X1 port map( A1 => n14928, A2 => n15080, B1 => n9141, B2 => 
                           n14926, ZN => n1860);
   U12267 : OAI22_X1 port map( A1 => n14928, A2 => n15083, B1 => n9140, B2 => 
                           n14926, ZN => n1861);
   U12268 : OAI22_X1 port map( A1 => n14928, A2 => n15086, B1 => n9139, B2 => 
                           n14926, ZN => n1862);
   U12269 : OAI22_X1 port map( A1 => n14928, A2 => n15089, B1 => n9138, B2 => 
                           n14926, ZN => n1863);
   U12270 : OAI22_X1 port map( A1 => n14929, A2 => n15092, B1 => n9137, B2 => 
                           n14926, ZN => n1864);
   U12271 : OAI22_X1 port map( A1 => n14929, A2 => n15095, B1 => n9136, B2 => 
                           n14926, ZN => n1865);
   U12272 : OAI22_X1 port map( A1 => n14929, A2 => n15098, B1 => n9135, B2 => 
                           n12004, ZN => n1866);
   U12273 : OAI22_X1 port map( A1 => n14929, A2 => n15101, B1 => n9134, B2 => 
                           n12004, ZN => n1867);
   U12274 : OAI22_X1 port map( A1 => n14929, A2 => n15104, B1 => n9133, B2 => 
                           n12004, ZN => n1868);
   U12275 : OAI22_X1 port map( A1 => n14930, A2 => n15107, B1 => n9132, B2 => 
                           n14926, ZN => n1869);
   U12276 : OAI22_X1 port map( A1 => n14930, A2 => n15110, B1 => n9131, B2 => 
                           n14926, ZN => n1870);
   U12277 : OAI22_X1 port map( A1 => n14930, A2 => n15113, B1 => n9130, B2 => 
                           n14926, ZN => n1871);
   U12278 : OAI22_X1 port map( A1 => n14930, A2 => n15116, B1 => n9129, B2 => 
                           n14926, ZN => n1872);
   U12279 : OAI22_X1 port map( A1 => n14930, A2 => n15119, B1 => n9128, B2 => 
                           n14926, ZN => n1873);
   U12280 : OAI22_X1 port map( A1 => n14931, A2 => n15122, B1 => n9127, B2 => 
                           n14926, ZN => n1874);
   U12281 : OAI22_X1 port map( A1 => n14931, A2 => n15125, B1 => n9126, B2 => 
                           n14926, ZN => n1875);
   U12282 : OAI22_X1 port map( A1 => n14931, A2 => n15128, B1 => n9125, B2 => 
                           n14926, ZN => n1876);
   U12283 : OAI22_X1 port map( A1 => n14931, A2 => n15131, B1 => n9124, B2 => 
                           n14926, ZN => n1877);
   U12284 : OAI22_X1 port map( A1 => n14963, A2 => n15061, B1 => n9019, B2 => 
                           n14962, ZN => n1982);
   U12285 : OAI22_X1 port map( A1 => n14963, A2 => n15064, B1 => n9018, B2 => 
                           n14962, ZN => n1983);
   U12286 : OAI22_X1 port map( A1 => n14963, A2 => n15067, B1 => n9017, B2 => 
                           n14962, ZN => n1984);
   U12287 : OAI22_X1 port map( A1 => n14963, A2 => n15070, B1 => n9016, B2 => 
                           n14962, ZN => n1985);
   U12288 : OAI22_X1 port map( A1 => n14963, A2 => n15073, B1 => n9015, B2 => 
                           n14962, ZN => n1986);
   U12289 : OAI22_X1 port map( A1 => n14964, A2 => n15076, B1 => n9014, B2 => 
                           n14962, ZN => n1987);
   U12290 : OAI22_X1 port map( A1 => n14964, A2 => n15079, B1 => n9013, B2 => 
                           n14962, ZN => n1988);
   U12291 : OAI22_X1 port map( A1 => n14964, A2 => n15082, B1 => n9012, B2 => 
                           n14962, ZN => n1989);
   U12292 : OAI22_X1 port map( A1 => n14964, A2 => n15085, B1 => n9011, B2 => 
                           n14962, ZN => n1990);
   U12293 : OAI22_X1 port map( A1 => n14964, A2 => n15088, B1 => n9010, B2 => 
                           n14962, ZN => n1991);
   U12294 : OAI22_X1 port map( A1 => n14965, A2 => n15091, B1 => n9009, B2 => 
                           n14962, ZN => n1992);
   U12295 : OAI22_X1 port map( A1 => n14965, A2 => n15094, B1 => n9008, B2 => 
                           n14962, ZN => n1993);
   U12296 : OAI22_X1 port map( A1 => n14965, A2 => n15097, B1 => n9007, B2 => 
                           n11999, ZN => n1994);
   U12297 : OAI22_X1 port map( A1 => n14965, A2 => n15100, B1 => n9006, B2 => 
                           n11999, ZN => n1995);
   U12298 : OAI22_X1 port map( A1 => n14965, A2 => n15103, B1 => n9005, B2 => 
                           n11999, ZN => n1996);
   U12299 : OAI22_X1 port map( A1 => n14966, A2 => n15106, B1 => n9004, B2 => 
                           n14962, ZN => n1997);
   U12300 : OAI22_X1 port map( A1 => n14966, A2 => n15109, B1 => n9003, B2 => 
                           n14962, ZN => n1998);
   U12301 : OAI22_X1 port map( A1 => n14966, A2 => n15112, B1 => n9002, B2 => 
                           n14962, ZN => n1999);
   U12302 : OAI22_X1 port map( A1 => n14966, A2 => n15115, B1 => n9001, B2 => 
                           n14962, ZN => n2000);
   U12303 : OAI22_X1 port map( A1 => n14966, A2 => n15118, B1 => n9000, B2 => 
                           n14962, ZN => n2001);
   U12304 : OAI22_X1 port map( A1 => n14967, A2 => n15121, B1 => n8999, B2 => 
                           n14962, ZN => n2002);
   U12305 : OAI22_X1 port map( A1 => n14967, A2 => n15124, B1 => n8998, B2 => 
                           n14962, ZN => n2003);
   U12306 : OAI22_X1 port map( A1 => n14967, A2 => n15127, B1 => n8997, B2 => 
                           n14962, ZN => n2004);
   U12307 : OAI22_X1 port map( A1 => n14967, A2 => n15130, B1 => n8996, B2 => 
                           n14962, ZN => n2005);
   U12308 : OAI221_X1 port map( B1 => n13824, B2 => n14681, C1 => n13216, C2 =>
                           n14676, A => n12768, ZN => n12767);
   U12309 : OAI21_X1 port map( B1 => n12769, B2 => n12770, A => n14675, ZN => 
                           n12768);
   U12310 : OAI221_X1 port map( B1 => n9635, B2 => n14662, C1 => n13892, C2 => 
                           n14659, A => n12772, ZN => n12769);
   U12311 : OAI221_X1 port map( B1 => n9507, B2 => n14671, C1 => n13893, C2 => 
                           n14669, A => n12771, ZN => n12770);
   U12312 : OAI221_X1 port map( B1 => n13825, B2 => n14681, C1 => n13217, C2 =>
                           n14676, A => n12751, ZN => n12750);
   U12313 : OAI21_X1 port map( B1 => n12752, B2 => n12753, A => n14675, ZN => 
                           n12751);
   U12314 : OAI221_X1 port map( B1 => n9634, B2 => n14662, C1 => n13894, C2 => 
                           n14660, A => n12755, ZN => n12752);
   U12315 : OAI221_X1 port map( B1 => n9506, B2 => n14672, C1 => n13895, C2 => 
                           n14670, A => n12754, ZN => n12753);
   U12316 : OAI221_X1 port map( B1 => n13826, B2 => n14681, C1 => n13218, C2 =>
                           n14676, A => n12734, ZN => n12733);
   U12317 : OAI21_X1 port map( B1 => n12735, B2 => n12736, A => n14675, ZN => 
                           n12734);
   U12318 : OAI221_X1 port map( B1 => n9633, B2 => n14662, C1 => n13896, C2 => 
                           n14659, A => n12738, ZN => n12735);
   U12319 : OAI221_X1 port map( B1 => n9505, B2 => n14671, C1 => n13897, C2 => 
                           n14669, A => n12737, ZN => n12736);
   U12320 : OAI221_X1 port map( B1 => n13827, B2 => n14681, C1 => n13219, C2 =>
                           n14676, A => n12717, ZN => n12716);
   U12321 : OAI21_X1 port map( B1 => n12718, B2 => n12719, A => n14675, ZN => 
                           n12717);
   U12322 : OAI221_X1 port map( B1 => n9632, B2 => n14662, C1 => n13898, C2 => 
                           n14660, A => n12721, ZN => n12718);
   U12323 : OAI221_X1 port map( B1 => n9504, B2 => n14672, C1 => n13899, C2 => 
                           n14670, A => n12720, ZN => n12719);
   U12324 : OAI221_X1 port map( B1 => n13828, B2 => n14681, C1 => n13220, C2 =>
                           n14676, A => n12700, ZN => n12699);
   U12325 : OAI21_X1 port map( B1 => n12701, B2 => n12702, A => n14675, ZN => 
                           n12700);
   U12326 : OAI221_X1 port map( B1 => n9631, B2 => n14662, C1 => n13900, C2 => 
                           n14659, A => n12704, ZN => n12701);
   U12327 : OAI221_X1 port map( B1 => n9503, B2 => n14671, C1 => n13901, C2 => 
                           n14669, A => n12703, ZN => n12702);
   U12328 : OAI221_X1 port map( B1 => n13829, B2 => n14681, C1 => n13221, C2 =>
                           n14676, A => n12683, ZN => n12682);
   U12329 : OAI21_X1 port map( B1 => n12684, B2 => n12685, A => n14675, ZN => 
                           n12683);
   U12330 : OAI221_X1 port map( B1 => n9630, B2 => n14662, C1 => n13902, C2 => 
                           n14660, A => n12687, ZN => n12684);
   U12331 : OAI221_X1 port map( B1 => n9502, B2 => n14672, C1 => n13903, C2 => 
                           n14670, A => n12686, ZN => n12685);
   U12332 : OAI221_X1 port map( B1 => n13830, B2 => n14681, C1 => n13188, C2 =>
                           n14676, A => n12666, ZN => n12665);
   U12333 : OAI21_X1 port map( B1 => n12667, B2 => n12668, A => n14675, ZN => 
                           n12666);
   U12334 : OAI221_X1 port map( B1 => n13636, B2 => n14662, C1 => n13904, C2 =>
                           n14659, A => n12670, ZN => n12667);
   U12335 : OAI221_X1 port map( B1 => n9501, B2 => n14671, C1 => n13905, C2 => 
                           n14669, A => n12669, ZN => n12668);
   U12336 : OAI221_X1 port map( B1 => n13831, B2 => n14681, C1 => n13189, C2 =>
                           n14677, A => n12617, ZN => n12614);
   U12337 : OAI21_X1 port map( B1 => n12618, B2 => n12619, A => n14675, ZN => 
                           n12617);
   U12338 : OAI221_X1 port map( B1 => n13727, B2 => n14662, C1 => n13906, C2 =>
                           n14660, A => n12628, ZN => n12618);
   U12339 : OAI221_X1 port map( B1 => n9500, B2 => n14672, C1 => n13907, C2 => 
                           n14670, A => n12623, ZN => n12619);
   U12340 : OAI221_X1 port map( B1 => n13824, B2 => n14779, C1 => n13246, C2 =>
                           n14774, A => n12187, ZN => n12186);
   U12341 : OAI21_X1 port map( B1 => n12188, B2 => n12189, A => n14773, ZN => 
                           n12187);
   U12342 : OAI221_X1 port map( B1 => n9635, B2 => n14760, C1 => n13892, C2 => 
                           n14757, A => n12191, ZN => n12188);
   U12343 : OAI221_X1 port map( B1 => n9507, B2 => n14769, C1 => n13893, C2 => 
                           n14767, A => n12190, ZN => n12189);
   U12344 : OAI221_X1 port map( B1 => n13825, B2 => n14779, C1 => n13247, C2 =>
                           n14774, A => n12170, ZN => n12169);
   U12345 : OAI21_X1 port map( B1 => n12171, B2 => n12172, A => n14773, ZN => 
                           n12170);
   U12346 : OAI221_X1 port map( B1 => n9634, B2 => n14760, C1 => n13894, C2 => 
                           n14758, A => n12174, ZN => n12171);
   U12347 : OAI221_X1 port map( B1 => n9506, B2 => n14770, C1 => n13895, C2 => 
                           n14768, A => n12173, ZN => n12172);
   U12348 : OAI221_X1 port map( B1 => n13826, B2 => n14779, C1 => n13248, C2 =>
                           n14774, A => n12153, ZN => n12152);
   U12349 : OAI21_X1 port map( B1 => n12154, B2 => n12155, A => n14773, ZN => 
                           n12153);
   U12350 : OAI221_X1 port map( B1 => n9633, B2 => n14760, C1 => n13896, C2 => 
                           n14757, A => n12157, ZN => n12154);
   U12351 : OAI221_X1 port map( B1 => n9505, B2 => n14769, C1 => n13897, C2 => 
                           n14767, A => n12156, ZN => n12155);
   U12352 : OAI221_X1 port map( B1 => n13827, B2 => n14779, C1 => n13249, C2 =>
                           n14774, A => n12136, ZN => n12135);
   U12353 : OAI21_X1 port map( B1 => n12137, B2 => n12138, A => n14773, ZN => 
                           n12136);
   U12354 : OAI221_X1 port map( B1 => n9632, B2 => n14760, C1 => n13898, C2 => 
                           n14758, A => n12140, ZN => n12137);
   U12355 : OAI221_X1 port map( B1 => n9504, B2 => n14770, C1 => n13899, C2 => 
                           n14768, A => n12139, ZN => n12138);
   U12356 : OAI221_X1 port map( B1 => n13828, B2 => n14779, C1 => n13250, C2 =>
                           n14774, A => n12119, ZN => n12118);
   U12357 : OAI21_X1 port map( B1 => n12120, B2 => n12121, A => n14773, ZN => 
                           n12119);
   U12358 : OAI221_X1 port map( B1 => n9631, B2 => n14760, C1 => n13900, C2 => 
                           n14757, A => n12123, ZN => n12120);
   U12359 : OAI221_X1 port map( B1 => n9503, B2 => n14769, C1 => n13901, C2 => 
                           n14767, A => n12122, ZN => n12121);
   U12360 : OAI221_X1 port map( B1 => n13829, B2 => n14779, C1 => n13251, C2 =>
                           n14774, A => n12102, ZN => n12101);
   U12361 : OAI21_X1 port map( B1 => n12103, B2 => n12104, A => n14773, ZN => 
                           n12102);
   U12362 : OAI221_X1 port map( B1 => n9630, B2 => n14760, C1 => n13902, C2 => 
                           n14758, A => n12106, ZN => n12103);
   U12363 : OAI221_X1 port map( B1 => n9502, B2 => n14770, C1 => n13903, C2 => 
                           n14768, A => n12105, ZN => n12104);
   U12364 : OAI221_X1 port map( B1 => n13830, B2 => n14779, C1 => n13190, C2 =>
                           n14774, A => n12085, ZN => n12084);
   U12365 : OAI21_X1 port map( B1 => n12086, B2 => n12087, A => n14773, ZN => 
                           n12085);
   U12366 : OAI221_X1 port map( B1 => n13636, B2 => n14760, C1 => n13904, C2 =>
                           n14757, A => n12089, ZN => n12086);
   U12367 : OAI221_X1 port map( B1 => n9501, B2 => n14769, C1 => n13905, C2 => 
                           n14767, A => n12088, ZN => n12087);
   U12368 : OAI221_X1 port map( B1 => n13831, B2 => n14779, C1 => n13191, C2 =>
                           n14775, A => n12036, ZN => n12033);
   U12369 : OAI21_X1 port map( B1 => n12037, B2 => n12038, A => n14773, ZN => 
                           n12036);
   U12370 : OAI221_X1 port map( B1 => n13727, B2 => n14760, C1 => n13906, C2 =>
                           n14758, A => n12047, ZN => n12037);
   U12371 : OAI221_X1 port map( B1 => n9500, B2 => n14770, C1 => n13907, C2 => 
                           n14768, A => n12042, ZN => n12038);
   U12372 : OAI221_X1 port map( B1 => n14086, B2 => n14679, C1 => n13192, C2 =>
                           n14678, A => n13176, ZN => n13175);
   U12373 : OAI21_X1 port map( B1 => n13177, B2 => n13178, A => n14673, ZN => 
                           n13176);
   U12374 : OAI221_X1 port map( B1 => n9659, B2 => n14661, C1 => n13908, C2 => 
                           n14659, A => n13180, ZN => n13177);
   U12375 : OAI221_X1 port map( B1 => n9531, B2 => n14671, C1 => n14218, C2 => 
                           n14669, A => n13179, ZN => n13178);
   U12376 : OAI221_X1 port map( B1 => n14087, B2 => n14679, C1 => n13193, C2 =>
                           n14678, A => n13159, ZN => n13158);
   U12377 : OAI21_X1 port map( B1 => n13160, B2 => n13161, A => n14673, ZN => 
                           n13159);
   U12378 : OAI221_X1 port map( B1 => n13637, B2 => n14662, C1 => n13909, C2 =>
                           n14659, A => n13163, ZN => n13160);
   U12379 : OAI221_X1 port map( B1 => n9530, B2 => n14671, C1 => n14219, C2 => 
                           n14669, A => n13162, ZN => n13161);
   U12380 : OAI221_X1 port map( B1 => n14088, B2 => n14679, C1 => n13194, C2 =>
                           n14678, A => n13142, ZN => n13141);
   U12381 : OAI21_X1 port map( B1 => n13143, B2 => n13144, A => n14673, ZN => 
                           n13142);
   U12382 : OAI221_X1 port map( B1 => n13638, B2 => n14661, C1 => n13910, C2 =>
                           n14659, A => n13146, ZN => n13143);
   U12383 : OAI221_X1 port map( B1 => n9529, B2 => n14671, C1 => n14220, C2 => 
                           n14669, A => n13145, ZN => n13144);
   U12384 : OAI221_X1 port map( B1 => n14089, B2 => n14679, C1 => n13195, C2 =>
                           n14678, A => n13125, ZN => n13124);
   U12385 : OAI21_X1 port map( B1 => n13126, B2 => n13127, A => n14673, ZN => 
                           n13125);
   U12386 : OAI221_X1 port map( B1 => n13639, B2 => n14662, C1 => n13911, C2 =>
                           n14659, A => n13129, ZN => n13126);
   U12387 : OAI221_X1 port map( B1 => n9528, B2 => n14671, C1 => n14221, C2 => 
                           n14669, A => n13128, ZN => n13127);
   U12388 : OAI221_X1 port map( B1 => n14090, B2 => n14679, C1 => n13196, C2 =>
                           n14678, A => n13108, ZN => n13107);
   U12389 : OAI21_X1 port map( B1 => n13109, B2 => n13110, A => n14673, ZN => 
                           n13108);
   U12390 : OAI221_X1 port map( B1 => n13640, B2 => n14661, C1 => n13912, C2 =>
                           n14659, A => n13112, ZN => n13109);
   U12391 : OAI221_X1 port map( B1 => n9527, B2 => n14671, C1 => n14222, C2 => 
                           n14669, A => n13111, ZN => n13110);
   U12392 : OAI221_X1 port map( B1 => n14091, B2 => n14679, C1 => n13197, C2 =>
                           n14678, A => n13091, ZN => n13090);
   U12393 : OAI21_X1 port map( B1 => n13092, B2 => n13093, A => n14673, ZN => 
                           n13091);
   U12394 : OAI221_X1 port map( B1 => n13641, B2 => n14662, C1 => n13913, C2 =>
                           n14659, A => n13095, ZN => n13092);
   U12395 : OAI221_X1 port map( B1 => n9526, B2 => n14671, C1 => n14223, C2 => 
                           n14669, A => n13094, ZN => n13093);
   U12396 : OAI221_X1 port map( B1 => n14092, B2 => n14679, C1 => n13198, C2 =>
                           n14678, A => n13074, ZN => n13073);
   U12397 : OAI21_X1 port map( B1 => n13075, B2 => n13076, A => n14673, ZN => 
                           n13074);
   U12398 : OAI221_X1 port map( B1 => n13642, B2 => n14661, C1 => n13914, C2 =>
                           n14659, A => n13078, ZN => n13075);
   U12399 : OAI221_X1 port map( B1 => n9525, B2 => n14671, C1 => n14224, C2 => 
                           n14669, A => n13077, ZN => n13076);
   U12400 : OAI221_X1 port map( B1 => n14093, B2 => n14679, C1 => n13199, C2 =>
                           n14678, A => n13057, ZN => n13056);
   U12401 : OAI21_X1 port map( B1 => n13058, B2 => n13059, A => n14673, ZN => 
                           n13057);
   U12402 : OAI221_X1 port map( B1 => n13643, B2 => n14662, C1 => n13915, C2 =>
                           n14659, A => n13061, ZN => n13058);
   U12403 : OAI221_X1 port map( B1 => n9524, B2 => n14671, C1 => n14225, C2 => 
                           n14669, A => n13060, ZN => n13059);
   U12404 : OAI221_X1 port map( B1 => n14086, B2 => n14777, C1 => n13222, C2 =>
                           n14776, A => n12595, ZN => n12594);
   U12405 : OAI21_X1 port map( B1 => n12596, B2 => n12597, A => n14771, ZN => 
                           n12595);
   U12406 : OAI221_X1 port map( B1 => n9659, B2 => n14759, C1 => n13908, C2 => 
                           n14757, A => n12599, ZN => n12596);
   U12407 : OAI221_X1 port map( B1 => n9531, B2 => n14769, C1 => n14218, C2 => 
                           n14767, A => n12598, ZN => n12597);
   U12408 : OAI221_X1 port map( B1 => n14087, B2 => n14777, C1 => n13223, C2 =>
                           n14776, A => n12578, ZN => n12577);
   U12409 : OAI21_X1 port map( B1 => n12579, B2 => n12580, A => n14771, ZN => 
                           n12578);
   U12410 : OAI221_X1 port map( B1 => n13637, B2 => n14760, C1 => n13909, C2 =>
                           n14757, A => n12582, ZN => n12579);
   U12411 : OAI221_X1 port map( B1 => n9530, B2 => n14769, C1 => n14219, C2 => 
                           n14767, A => n12581, ZN => n12580);
   U12412 : OAI221_X1 port map( B1 => n14088, B2 => n14777, C1 => n13224, C2 =>
                           n14776, A => n12561, ZN => n12560);
   U12413 : OAI21_X1 port map( B1 => n12562, B2 => n12563, A => n14771, ZN => 
                           n12561);
   U12414 : OAI221_X1 port map( B1 => n13638, B2 => n14759, C1 => n13910, C2 =>
                           n14757, A => n12565, ZN => n12562);
   U12415 : OAI221_X1 port map( B1 => n9529, B2 => n14769, C1 => n14220, C2 => 
                           n14767, A => n12564, ZN => n12563);
   U12416 : OAI221_X1 port map( B1 => n14089, B2 => n14777, C1 => n13225, C2 =>
                           n14776, A => n12544, ZN => n12543);
   U12417 : OAI21_X1 port map( B1 => n12545, B2 => n12546, A => n14771, ZN => 
                           n12544);
   U12418 : OAI221_X1 port map( B1 => n13639, B2 => n14760, C1 => n13911, C2 =>
                           n14757, A => n12548, ZN => n12545);
   U12419 : OAI221_X1 port map( B1 => n9528, B2 => n14769, C1 => n14221, C2 => 
                           n14767, A => n12547, ZN => n12546);
   U12420 : OAI221_X1 port map( B1 => n14090, B2 => n14777, C1 => n13226, C2 =>
                           n14776, A => n12527, ZN => n12526);
   U12421 : OAI21_X1 port map( B1 => n12528, B2 => n12529, A => n14771, ZN => 
                           n12527);
   U12422 : OAI221_X1 port map( B1 => n13640, B2 => n14759, C1 => n13912, C2 =>
                           n14757, A => n12531, ZN => n12528);
   U12423 : OAI221_X1 port map( B1 => n9527, B2 => n14769, C1 => n14222, C2 => 
                           n14767, A => n12530, ZN => n12529);
   U12424 : OAI221_X1 port map( B1 => n14091, B2 => n14777, C1 => n13227, C2 =>
                           n14776, A => n12510, ZN => n12509);
   U12425 : OAI21_X1 port map( B1 => n12511, B2 => n12512, A => n14771, ZN => 
                           n12510);
   U12426 : OAI221_X1 port map( B1 => n13641, B2 => n14760, C1 => n13913, C2 =>
                           n14757, A => n12514, ZN => n12511);
   U12427 : OAI221_X1 port map( B1 => n9526, B2 => n14769, C1 => n14223, C2 => 
                           n14767, A => n12513, ZN => n12512);
   U12428 : OAI221_X1 port map( B1 => n14092, B2 => n14777, C1 => n13228, C2 =>
                           n14776, A => n12493, ZN => n12492);
   U12429 : OAI21_X1 port map( B1 => n12494, B2 => n12495, A => n14771, ZN => 
                           n12493);
   U12430 : OAI221_X1 port map( B1 => n13642, B2 => n14759, C1 => n13914, C2 =>
                           n14757, A => n12497, ZN => n12494);
   U12431 : OAI221_X1 port map( B1 => n9525, B2 => n14769, C1 => n14224, C2 => 
                           n14767, A => n12496, ZN => n12495);
   U12432 : OAI221_X1 port map( B1 => n14093, B2 => n14777, C1 => n13229, C2 =>
                           n14776, A => n12476, ZN => n12475);
   U12433 : OAI21_X1 port map( B1 => n12477, B2 => n12478, A => n14771, ZN => 
                           n12476);
   U12434 : OAI221_X1 port map( B1 => n13643, B2 => n14760, C1 => n13915, C2 =>
                           n14757, A => n12480, ZN => n12477);
   U12435 : OAI221_X1 port map( B1 => n9524, B2 => n14769, C1 => n14225, C2 => 
                           n14767, A => n12479, ZN => n12478);
   U12436 : NAND4_X1 port map( A1 => n13168, A2 => n13169, A3 => n13170, A4 => 
                           n13171, ZN => n1278);
   U12437 : AOI222_X1 port map( A1 => n14590, A2 => n14226, B1 => n14589, B2 =>
                           n13396, C1 => n14586, C2 => n13348, ZN => n13168);
   U12438 : AOI222_X1 port map( A1 => n14599, A2 => n13372, B1 => n14598, B2 =>
                           n13540, C1 => n14595, C2 => n13492, ZN => n13169);
   U12439 : AOI211_X1 port map( C1 => n14620, C2 => n13516, A => n13185, B => 
                           n13186, ZN => n13170);
   U12440 : NAND4_X1 port map( A1 => n13151, A2 => n13152, A3 => n13153, A4 => 
                           n13154, ZN => n1279);
   U12441 : AOI222_X1 port map( A1 => n14590, A2 => n14227, B1 => n14589, B2 =>
                           n13397, C1 => n14586, C2 => n13349, ZN => n13151);
   U12442 : AOI222_X1 port map( A1 => n14599, A2 => n13373, B1 => n14598, B2 =>
                           n13541, C1 => n14595, C2 => n13493, ZN => n13152);
   U12443 : AOI211_X1 port map( C1 => n14620, C2 => n13517, A => n13165, B => 
                           n13166, ZN => n13153);
   U12444 : NAND4_X1 port map( A1 => n13134, A2 => n13135, A3 => n13136, A4 => 
                           n13137, ZN => n1280);
   U12445 : AOI222_X1 port map( A1 => n14590, A2 => n14228, B1 => n14589, B2 =>
                           n13398, C1 => n14586, C2 => n13350, ZN => n13134);
   U12446 : AOI222_X1 port map( A1 => n14599, A2 => n13374, B1 => n14598, B2 =>
                           n13542, C1 => n14595, C2 => n13494, ZN => n13135);
   U12447 : AOI211_X1 port map( C1 => n14620, C2 => n13518, A => n13148, B => 
                           n13149, ZN => n13136);
   U12448 : NAND4_X1 port map( A1 => n13117, A2 => n13118, A3 => n13119, A4 => 
                           n13120, ZN => n1281);
   U12449 : AOI222_X1 port map( A1 => n14590, A2 => n14229, B1 => n14589, B2 =>
                           n13399, C1 => n14586, C2 => n13351, ZN => n13117);
   U12450 : AOI222_X1 port map( A1 => n14599, A2 => n13375, B1 => n14598, B2 =>
                           n13543, C1 => n14595, C2 => n13495, ZN => n13118);
   U12451 : AOI211_X1 port map( C1 => n14620, C2 => n13519, A => n13131, B => 
                           n13132, ZN => n13119);
   U12452 : NAND4_X1 port map( A1 => n13100, A2 => n13101, A3 => n13102, A4 => 
                           n13103, ZN => n1282);
   U12453 : AOI222_X1 port map( A1 => n14590, A2 => n14230, B1 => n14589, B2 =>
                           n13400, C1 => n14586, C2 => n13352, ZN => n13100);
   U12454 : AOI222_X1 port map( A1 => n14599, A2 => n13376, B1 => n14598, B2 =>
                           n13544, C1 => n14595, C2 => n13496, ZN => n13101);
   U12455 : AOI211_X1 port map( C1 => n14620, C2 => n13520, A => n13114, B => 
                           n13115, ZN => n13102);
   U12456 : NAND4_X1 port map( A1 => n13083, A2 => n13084, A3 => n13085, A4 => 
                           n13086, ZN => n1283);
   U12457 : AOI222_X1 port map( A1 => n14590, A2 => n14231, B1 => n14589, B2 =>
                           n13401, C1 => n14586, C2 => n13353, ZN => n13083);
   U12458 : AOI222_X1 port map( A1 => n14599, A2 => n13377, B1 => n14598, B2 =>
                           n13545, C1 => n14595, C2 => n13497, ZN => n13084);
   U12459 : AOI211_X1 port map( C1 => n14620, C2 => n13521, A => n13097, B => 
                           n13098, ZN => n13085);
   U12460 : NAND4_X1 port map( A1 => n13066, A2 => n13067, A3 => n13068, A4 => 
                           n13069, ZN => n1284);
   U12461 : AOI222_X1 port map( A1 => n14590, A2 => n14232, B1 => n14589, B2 =>
                           n13402, C1 => n14586, C2 => n13354, ZN => n13066);
   U12462 : AOI222_X1 port map( A1 => n14599, A2 => n13378, B1 => n14598, B2 =>
                           n13546, C1 => n14595, C2 => n13498, ZN => n13067);
   U12463 : AOI211_X1 port map( C1 => n14620, C2 => n13522, A => n13080, B => 
                           n13081, ZN => n13068);
   U12464 : NAND4_X1 port map( A1 => n13049, A2 => n13050, A3 => n13051, A4 => 
                           n13052, ZN => n1285);
   U12465 : AOI222_X1 port map( A1 => n14590, A2 => n14233, B1 => n14589, B2 =>
                           n13403, C1 => n14586, C2 => n13355, ZN => n13049);
   U12466 : AOI222_X1 port map( A1 => n14599, A2 => n13379, B1 => n14598, B2 =>
                           n13547, C1 => n14595, C2 => n13499, ZN => n13050);
   U12467 : AOI211_X1 port map( C1 => n14620, C2 => n13523, A => n13063, B => 
                           n13064, ZN => n13051);
   U12468 : NAND4_X1 port map( A1 => n13032, A2 => n13033, A3 => n13034, A4 => 
                           n13035, ZN => n1286);
   U12469 : AOI222_X1 port map( A1 => n14590, A2 => n14234, B1 => n14588, B2 =>
                           n13404, C1 => n14585, C2 => n13356, ZN => n13032);
   U12470 : AOI222_X1 port map( A1 => n14599, A2 => n13380, B1 => n14597, B2 =>
                           n13548, C1 => n14594, C2 => n13500, ZN => n13033);
   U12471 : AOI211_X1 port map( C1 => n14620, C2 => n13524, A => n13046, B => 
                           n13047, ZN => n13034);
   U12472 : NAND4_X1 port map( A1 => n13015, A2 => n13016, A3 => n13017, A4 => 
                           n13018, ZN => n1287);
   U12473 : AOI222_X1 port map( A1 => n14590, A2 => n14235, B1 => n14588, B2 =>
                           n13405, C1 => n14585, C2 => n13357, ZN => n13015);
   U12474 : AOI222_X1 port map( A1 => n14599, A2 => n13381, B1 => n14597, B2 =>
                           n13549, C1 => n14594, C2 => n13501, ZN => n13016);
   U12475 : AOI211_X1 port map( C1 => n14620, C2 => n13525, A => n13029, B => 
                           n13030, ZN => n13017);
   U12476 : NAND4_X1 port map( A1 => n12998, A2 => n12999, A3 => n13000, A4 => 
                           n13001, ZN => n1288);
   U12477 : AOI222_X1 port map( A1 => n14590, A2 => n14236, B1 => n14588, B2 =>
                           n13406, C1 => n14585, C2 => n13358, ZN => n12998);
   U12478 : AOI222_X1 port map( A1 => n14599, A2 => n13382, B1 => n14597, B2 =>
                           n13550, C1 => n14594, C2 => n13502, ZN => n12999);
   U12479 : AOI211_X1 port map( C1 => n14620, C2 => n13526, A => n13012, B => 
                           n13013, ZN => n13000);
   U12480 : NAND4_X1 port map( A1 => n12981, A2 => n12982, A3 => n12983, A4 => 
                           n12984, ZN => n1289);
   U12481 : AOI222_X1 port map( A1 => n14590, A2 => n14237, B1 => n14588, B2 =>
                           n13407, C1 => n14585, C2 => n13359, ZN => n12981);
   U12482 : AOI222_X1 port map( A1 => n14599, A2 => n13383, B1 => n14597, B2 =>
                           n13551, C1 => n14594, C2 => n13503, ZN => n12982);
   U12483 : AOI211_X1 port map( C1 => n14620, C2 => n13527, A => n12995, B => 
                           n12996, ZN => n12983);
   U12484 : NAND4_X1 port map( A1 => n12964, A2 => n12965, A3 => n12966, A4 => 
                           n12967, ZN => n1290);
   U12485 : AOI222_X1 port map( A1 => n14591, A2 => n14238, B1 => n14588, B2 =>
                           n13408, C1 => n14585, C2 => n13360, ZN => n12964);
   U12486 : AOI222_X1 port map( A1 => n14600, A2 => n13384, B1 => n14597, B2 =>
                           n13552, C1 => n14594, C2 => n13504, ZN => n12965);
   U12487 : AOI211_X1 port map( C1 => n14621, C2 => n13528, A => n12978, B => 
                           n12979, ZN => n12966);
   U12488 : NAND4_X1 port map( A1 => n12947, A2 => n12948, A3 => n12949, A4 => 
                           n12950, ZN => n1291);
   U12489 : AOI222_X1 port map( A1 => n14591, A2 => n14239, B1 => n14588, B2 =>
                           n13409, C1 => n14585, C2 => n13361, ZN => n12947);
   U12490 : AOI222_X1 port map( A1 => n14600, A2 => n13385, B1 => n14597, B2 =>
                           n13553, C1 => n14594, C2 => n13505, ZN => n12948);
   U12491 : AOI211_X1 port map( C1 => n14621, C2 => n13529, A => n12961, B => 
                           n12962, ZN => n12949);
   U12492 : NAND4_X1 port map( A1 => n12930, A2 => n12931, A3 => n12932, A4 => 
                           n12933, ZN => n1292);
   U12493 : AOI222_X1 port map( A1 => n14591, A2 => n14240, B1 => n14588, B2 =>
                           n13410, C1 => n14585, C2 => n13362, ZN => n12930);
   U12494 : AOI222_X1 port map( A1 => n14600, A2 => n13386, B1 => n14597, B2 =>
                           n13554, C1 => n14594, C2 => n13506, ZN => n12931);
   U12495 : AOI211_X1 port map( C1 => n14621, C2 => n13530, A => n12944, B => 
                           n12945, ZN => n12932);
   U12496 : NAND4_X1 port map( A1 => n12913, A2 => n12914, A3 => n12915, A4 => 
                           n12916, ZN => n1293);
   U12497 : AOI222_X1 port map( A1 => n14591, A2 => n14241, B1 => n14588, B2 =>
                           n13411, C1 => n14585, C2 => n13363, ZN => n12913);
   U12498 : AOI222_X1 port map( A1 => n14600, A2 => n13387, B1 => n14597, B2 =>
                           n13555, C1 => n14594, C2 => n13507, ZN => n12914);
   U12499 : AOI211_X1 port map( C1 => n14621, C2 => n13531, A => n12927, B => 
                           n12928, ZN => n12915);
   U12500 : NAND4_X1 port map( A1 => n12896, A2 => n12897, A3 => n12898, A4 => 
                           n12899, ZN => n1294);
   U12501 : AOI222_X1 port map( A1 => n14591, A2 => n14242, B1 => n14588, B2 =>
                           n13412, C1 => n14585, C2 => n13364, ZN => n12896);
   U12502 : AOI222_X1 port map( A1 => n14600, A2 => n13388, B1 => n14597, B2 =>
                           n13556, C1 => n14594, C2 => n13508, ZN => n12897);
   U12503 : AOI211_X1 port map( C1 => n14621, C2 => n13532, A => n12910, B => 
                           n12911, ZN => n12898);
   U12504 : NAND4_X1 port map( A1 => n12879, A2 => n12880, A3 => n12881, A4 => 
                           n12882, ZN => n1295);
   U12505 : AOI222_X1 port map( A1 => n14591, A2 => n14243, B1 => n14588, B2 =>
                           n13413, C1 => n14585, C2 => n13365, ZN => n12879);
   U12506 : AOI222_X1 port map( A1 => n14600, A2 => n13389, B1 => n14597, B2 =>
                           n13557, C1 => n14594, C2 => n13509, ZN => n12880);
   U12507 : AOI211_X1 port map( C1 => n14621, C2 => n13533, A => n12893, B => 
                           n12894, ZN => n12881);
   U12508 : NAND4_X1 port map( A1 => n12862, A2 => n12863, A3 => n12864, A4 => 
                           n12865, ZN => n1296);
   U12509 : AOI222_X1 port map( A1 => n14591, A2 => n14244, B1 => n14588, B2 =>
                           n13414, C1 => n14585, C2 => n13366, ZN => n12862);
   U12510 : AOI222_X1 port map( A1 => n14600, A2 => n13390, B1 => n14597, B2 =>
                           n13558, C1 => n14594, C2 => n13510, ZN => n12863);
   U12511 : AOI211_X1 port map( C1 => n14621, C2 => n13534, A => n12876, B => 
                           n12877, ZN => n12864);
   U12512 : NAND4_X1 port map( A1 => n12845, A2 => n12846, A3 => n12847, A4 => 
                           n12848, ZN => n1297);
   U12513 : AOI222_X1 port map( A1 => n14591, A2 => n14245, B1 => n14588, B2 =>
                           n13415, C1 => n14585, C2 => n13367, ZN => n12845);
   U12514 : AOI222_X1 port map( A1 => n14600, A2 => n13391, B1 => n14597, B2 =>
                           n13559, C1 => n14594, C2 => n13511, ZN => n12846);
   U12515 : AOI211_X1 port map( C1 => n14621, C2 => n13535, A => n12859, B => 
                           n12860, ZN => n12847);
   U12516 : NAND4_X1 port map( A1 => n12828, A2 => n12829, A3 => n12830, A4 => 
                           n12831, ZN => n1298);
   U12517 : AOI222_X1 port map( A1 => n14591, A2 => n14246, B1 => n14587, B2 =>
                           n13416, C1 => n14584, C2 => n13368, ZN => n12828);
   U12518 : AOI222_X1 port map( A1 => n14600, A2 => n13392, B1 => n14596, B2 =>
                           n13560, C1 => n14593, C2 => n13512, ZN => n12829);
   U12519 : AOI211_X1 port map( C1 => n14621, C2 => n13536, A => n12842, B => 
                           n12843, ZN => n12830);
   U12520 : NAND4_X1 port map( A1 => n12811, A2 => n12812, A3 => n12813, A4 => 
                           n12814, ZN => n1299);
   U12521 : AOI222_X1 port map( A1 => n14591, A2 => n14247, B1 => n14587, B2 =>
                           n13417, C1 => n14584, C2 => n13369, ZN => n12811);
   U12522 : AOI222_X1 port map( A1 => n14600, A2 => n13393, B1 => n14596, B2 =>
                           n13561, C1 => n14593, C2 => n13513, ZN => n12812);
   U12523 : AOI211_X1 port map( C1 => n14621, C2 => n13537, A => n12825, B => 
                           n12826, ZN => n12813);
   U12524 : NAND4_X1 port map( A1 => n12794, A2 => n12795, A3 => n12796, A4 => 
                           n12797, ZN => n1300);
   U12525 : AOI222_X1 port map( A1 => n14591, A2 => n14248, B1 => n14587, B2 =>
                           n13418, C1 => n14584, C2 => n13370, ZN => n12794);
   U12526 : AOI222_X1 port map( A1 => n14600, A2 => n13394, B1 => n14596, B2 =>
                           n13562, C1 => n14593, C2 => n13514, ZN => n12795);
   U12527 : AOI211_X1 port map( C1 => n14621, C2 => n13538, A => n12808, B => 
                           n12809, ZN => n12796);
   U12528 : NAND4_X1 port map( A1 => n12777, A2 => n12778, A3 => n12779, A4 => 
                           n12780, ZN => n1301);
   U12529 : AOI222_X1 port map( A1 => n14591, A2 => n14249, B1 => n14587, B2 =>
                           n13419, C1 => n14584, C2 => n13371, ZN => n12777);
   U12530 : AOI222_X1 port map( A1 => n14600, A2 => n13395, B1 => n14596, B2 =>
                           n13563, C1 => n14593, C2 => n13515, ZN => n12778);
   U12531 : AOI211_X1 port map( C1 => n14621, C2 => n13539, A => n12791, B => 
                           n12792, ZN => n12779);
   U12532 : NAND4_X1 port map( A1 => n12760, A2 => n12761, A3 => n12762, A4 => 
                           n12763, ZN => n1302);
   U12533 : AOI222_X1 port map( A1 => n14592, A2 => n14250, B1 => n14587, B2 =>
                           n13316, C1 => n14584, C2 => n13300, ZN => n12760);
   U12534 : AOI222_X1 port map( A1 => n14601, A2 => n13308, B1 => n14596, B2 =>
                           n13268, C1 => n14593, C2 => n13252, ZN => n12761);
   U12535 : AOI211_X1 port map( C1 => n14622, C2 => n13260, A => n12774, B => 
                           n12775, ZN => n12762);
   U12536 : NAND4_X1 port map( A1 => n12743, A2 => n12744, A3 => n12745, A4 => 
                           n12746, ZN => n1303);
   U12537 : AOI222_X1 port map( A1 => n14592, A2 => n14251, B1 => n14587, B2 =>
                           n13317, C1 => n14584, C2 => n13301, ZN => n12743);
   U12538 : AOI222_X1 port map( A1 => n14601, A2 => n13309, B1 => n14596, B2 =>
                           n13269, C1 => n14593, C2 => n13253, ZN => n12744);
   U12539 : AOI211_X1 port map( C1 => n14622, C2 => n13261, A => n12757, B => 
                           n12758, ZN => n12745);
   U12540 : NAND4_X1 port map( A1 => n12726, A2 => n12727, A3 => n12728, A4 => 
                           n12729, ZN => n1304);
   U12541 : AOI222_X1 port map( A1 => n14592, A2 => n14252, B1 => n14587, B2 =>
                           n13318, C1 => n14584, C2 => n13302, ZN => n12726);
   U12542 : AOI222_X1 port map( A1 => n14601, A2 => n13310, B1 => n14596, B2 =>
                           n13270, C1 => n14593, C2 => n13254, ZN => n12727);
   U12543 : AOI211_X1 port map( C1 => n14622, C2 => n13262, A => n12740, B => 
                           n12741, ZN => n12728);
   U12544 : NAND4_X1 port map( A1 => n12709, A2 => n12710, A3 => n12711, A4 => 
                           n12712, ZN => n1305);
   U12545 : AOI222_X1 port map( A1 => n14592, A2 => n14253, B1 => n14587, B2 =>
                           n13319, C1 => n14584, C2 => n13303, ZN => n12709);
   U12546 : AOI222_X1 port map( A1 => n14601, A2 => n13311, B1 => n14596, B2 =>
                           n13271, C1 => n14593, C2 => n13255, ZN => n12710);
   U12547 : AOI211_X1 port map( C1 => n14622, C2 => n13263, A => n12723, B => 
                           n12724, ZN => n12711);
   U12548 : NAND4_X1 port map( A1 => n12692, A2 => n12693, A3 => n12694, A4 => 
                           n12695, ZN => n1306);
   U12549 : AOI222_X1 port map( A1 => n14592, A2 => n14254, B1 => n14587, B2 =>
                           n13320, C1 => n14584, C2 => n13304, ZN => n12692);
   U12550 : AOI222_X1 port map( A1 => n14601, A2 => n13312, B1 => n14596, B2 =>
                           n13272, C1 => n14593, C2 => n13256, ZN => n12693);
   U12551 : AOI211_X1 port map( C1 => n14622, C2 => n13264, A => n12706, B => 
                           n12707, ZN => n12694);
   U12552 : NAND4_X1 port map( A1 => n12675, A2 => n12676, A3 => n12677, A4 => 
                           n12678, ZN => n1307);
   U12553 : AOI222_X1 port map( A1 => n14592, A2 => n14255, B1 => n14587, B2 =>
                           n13321, C1 => n14584, C2 => n13305, ZN => n12675);
   U12554 : AOI222_X1 port map( A1 => n14601, A2 => n13313, B1 => n14596, B2 =>
                           n13273, C1 => n14593, C2 => n13257, ZN => n12676);
   U12555 : AOI211_X1 port map( C1 => n14622, C2 => n13265, A => n12689, B => 
                           n12690, ZN => n12677);
   U12556 : NAND4_X1 port map( A1 => n12658, A2 => n12659, A3 => n12660, A4 => 
                           n12661, ZN => n1308);
   U12557 : AOI222_X1 port map( A1 => n14592, A2 => n14256, B1 => n14587, B2 =>
                           n13322, C1 => n14584, C2 => n13306, ZN => n12658);
   U12558 : AOI222_X1 port map( A1 => n14601, A2 => n13314, B1 => n14596, B2 =>
                           n13274, C1 => n14593, C2 => n13258, ZN => n12659);
   U12559 : AOI211_X1 port map( C1 => n14622, C2 => n13266, A => n12672, B => 
                           n12673, ZN => n12660);
   U12560 : NAND4_X1 port map( A1 => n12607, A2 => n12608, A3 => n12609, A4 => 
                           n12610, ZN => n1309);
   U12561 : AOI222_X1 port map( A1 => n14592, A2 => n14257, B1 => n14587, B2 =>
                           n13323, C1 => n14584, C2 => n13307, ZN => n12607);
   U12562 : AOI222_X1 port map( A1 => n14601, A2 => n13315, B1 => n14596, B2 =>
                           n13275, C1 => n14593, C2 => n13259, ZN => n12608);
   U12563 : AOI211_X1 port map( C1 => n14622, C2 => n13267, A => n12643, B => 
                           n12644, ZN => n12609);
   U12564 : NAND4_X1 port map( A1 => n12587, A2 => n12588, A3 => n12589, A4 => 
                           n12590, ZN => n1310);
   U12565 : AOI222_X1 port map( A1 => n14688, A2 => n14226, B1 => n14687, B2 =>
                           n13396, C1 => n14684, C2 => n13348, ZN => n12587);
   U12566 : AOI222_X1 port map( A1 => n14697, A2 => n13372, B1 => n14696, B2 =>
                           n13540, C1 => n14693, C2 => n13492, ZN => n12588);
   U12567 : AOI211_X1 port map( C1 => n14718, C2 => n13516, A => n12604, B => 
                           n12605, ZN => n12589);
   U12568 : NAND4_X1 port map( A1 => n12570, A2 => n12571, A3 => n12572, A4 => 
                           n12573, ZN => n1311);
   U12569 : AOI222_X1 port map( A1 => n14688, A2 => n14227, B1 => n14687, B2 =>
                           n13397, C1 => n14684, C2 => n13349, ZN => n12570);
   U12570 : AOI222_X1 port map( A1 => n14697, A2 => n13373, B1 => n14696, B2 =>
                           n13541, C1 => n14693, C2 => n13493, ZN => n12571);
   U12571 : AOI211_X1 port map( C1 => n14718, C2 => n13517, A => n12584, B => 
                           n12585, ZN => n12572);
   U12572 : NAND4_X1 port map( A1 => n12553, A2 => n12554, A3 => n12555, A4 => 
                           n12556, ZN => n1312);
   U12573 : AOI222_X1 port map( A1 => n14688, A2 => n14228, B1 => n14687, B2 =>
                           n13398, C1 => n14684, C2 => n13350, ZN => n12553);
   U12574 : AOI222_X1 port map( A1 => n14697, A2 => n13374, B1 => n14696, B2 =>
                           n13542, C1 => n14693, C2 => n13494, ZN => n12554);
   U12575 : AOI211_X1 port map( C1 => n14718, C2 => n13518, A => n12567, B => 
                           n12568, ZN => n12555);
   U12576 : NAND4_X1 port map( A1 => n12536, A2 => n12537, A3 => n12538, A4 => 
                           n12539, ZN => n1313);
   U12577 : AOI222_X1 port map( A1 => n14688, A2 => n14229, B1 => n14687, B2 =>
                           n13399, C1 => n14684, C2 => n13351, ZN => n12536);
   U12578 : AOI222_X1 port map( A1 => n14697, A2 => n13375, B1 => n14696, B2 =>
                           n13543, C1 => n14693, C2 => n13495, ZN => n12537);
   U12579 : AOI211_X1 port map( C1 => n14718, C2 => n13519, A => n12550, B => 
                           n12551, ZN => n12538);
   U12580 : NAND4_X1 port map( A1 => n12519, A2 => n12520, A3 => n12521, A4 => 
                           n12522, ZN => n1314);
   U12581 : AOI222_X1 port map( A1 => n14688, A2 => n14230, B1 => n14687, B2 =>
                           n13400, C1 => n14684, C2 => n13352, ZN => n12519);
   U12582 : AOI222_X1 port map( A1 => n14697, A2 => n13376, B1 => n14696, B2 =>
                           n13544, C1 => n14693, C2 => n13496, ZN => n12520);
   U12583 : AOI211_X1 port map( C1 => n14718, C2 => n13520, A => n12533, B => 
                           n12534, ZN => n12521);
   U12584 : NAND4_X1 port map( A1 => n12502, A2 => n12503, A3 => n12504, A4 => 
                           n12505, ZN => n1315);
   U12585 : AOI222_X1 port map( A1 => n14688, A2 => n14231, B1 => n14687, B2 =>
                           n13401, C1 => n14684, C2 => n13353, ZN => n12502);
   U12586 : AOI222_X1 port map( A1 => n14697, A2 => n13377, B1 => n14696, B2 =>
                           n13545, C1 => n14693, C2 => n13497, ZN => n12503);
   U12587 : AOI211_X1 port map( C1 => n14718, C2 => n13521, A => n12516, B => 
                           n12517, ZN => n12504);
   U12588 : NAND4_X1 port map( A1 => n12485, A2 => n12486, A3 => n12487, A4 => 
                           n12488, ZN => n1316);
   U12589 : AOI222_X1 port map( A1 => n14688, A2 => n14232, B1 => n14687, B2 =>
                           n13402, C1 => n14684, C2 => n13354, ZN => n12485);
   U12590 : AOI222_X1 port map( A1 => n14697, A2 => n13378, B1 => n14696, B2 =>
                           n13546, C1 => n14693, C2 => n13498, ZN => n12486);
   U12591 : AOI211_X1 port map( C1 => n14718, C2 => n13522, A => n12499, B => 
                           n12500, ZN => n12487);
   U12592 : NAND4_X1 port map( A1 => n12468, A2 => n12469, A3 => n12470, A4 => 
                           n12471, ZN => n1317);
   U12593 : AOI222_X1 port map( A1 => n14688, A2 => n14233, B1 => n14687, B2 =>
                           n13403, C1 => n14684, C2 => n13355, ZN => n12468);
   U12594 : AOI222_X1 port map( A1 => n14697, A2 => n13379, B1 => n14696, B2 =>
                           n13547, C1 => n14693, C2 => n13499, ZN => n12469);
   U12595 : AOI211_X1 port map( C1 => n14718, C2 => n13523, A => n12482, B => 
                           n12483, ZN => n12470);
   U12596 : NAND4_X1 port map( A1 => n12451, A2 => n12452, A3 => n12453, A4 => 
                           n12454, ZN => n1318);
   U12597 : AOI222_X1 port map( A1 => n14688, A2 => n14234, B1 => n14686, B2 =>
                           n13404, C1 => n14683, C2 => n13356, ZN => n12451);
   U12598 : AOI222_X1 port map( A1 => n14697, A2 => n13380, B1 => n14695, B2 =>
                           n13548, C1 => n14692, C2 => n13500, ZN => n12452);
   U12599 : AOI211_X1 port map( C1 => n14718, C2 => n13524, A => n12465, B => 
                           n12466, ZN => n12453);
   U12600 : NAND4_X1 port map( A1 => n12434, A2 => n12435, A3 => n12436, A4 => 
                           n12437, ZN => n1319);
   U12601 : AOI222_X1 port map( A1 => n14688, A2 => n14235, B1 => n14686, B2 =>
                           n13405, C1 => n14683, C2 => n13357, ZN => n12434);
   U12602 : AOI222_X1 port map( A1 => n14697, A2 => n13381, B1 => n14695, B2 =>
                           n13549, C1 => n14692, C2 => n13501, ZN => n12435);
   U12603 : AOI211_X1 port map( C1 => n14718, C2 => n13525, A => n12448, B => 
                           n12449, ZN => n12436);
   U12604 : NAND4_X1 port map( A1 => n12417, A2 => n12418, A3 => n12419, A4 => 
                           n12420, ZN => n1320);
   U12605 : AOI222_X1 port map( A1 => n14688, A2 => n14236, B1 => n14686, B2 =>
                           n13406, C1 => n14683, C2 => n13358, ZN => n12417);
   U12606 : AOI222_X1 port map( A1 => n14697, A2 => n13382, B1 => n14695, B2 =>
                           n13550, C1 => n14692, C2 => n13502, ZN => n12418);
   U12607 : AOI211_X1 port map( C1 => n14718, C2 => n13526, A => n12431, B => 
                           n12432, ZN => n12419);
   U12608 : NAND4_X1 port map( A1 => n12400, A2 => n12401, A3 => n12402, A4 => 
                           n12403, ZN => n1321);
   U12609 : AOI222_X1 port map( A1 => n14688, A2 => n14237, B1 => n14686, B2 =>
                           n13407, C1 => n14683, C2 => n13359, ZN => n12400);
   U12610 : AOI222_X1 port map( A1 => n14697, A2 => n13383, B1 => n14695, B2 =>
                           n13551, C1 => n14692, C2 => n13503, ZN => n12401);
   U12611 : AOI211_X1 port map( C1 => n14718, C2 => n13527, A => n12414, B => 
                           n12415, ZN => n12402);
   U12612 : NAND4_X1 port map( A1 => n12383, A2 => n12384, A3 => n12385, A4 => 
                           n12386, ZN => n1322);
   U12613 : AOI222_X1 port map( A1 => n14689, A2 => n14238, B1 => n14686, B2 =>
                           n13408, C1 => n14683, C2 => n13360, ZN => n12383);
   U12614 : AOI222_X1 port map( A1 => n14698, A2 => n13384, B1 => n14695, B2 =>
                           n13552, C1 => n14692, C2 => n13504, ZN => n12384);
   U12615 : AOI211_X1 port map( C1 => n14719, C2 => n13528, A => n12397, B => 
                           n12398, ZN => n12385);
   U12616 : NAND4_X1 port map( A1 => n12366, A2 => n12367, A3 => n12368, A4 => 
                           n12369, ZN => n1323);
   U12617 : AOI222_X1 port map( A1 => n14689, A2 => n14239, B1 => n14686, B2 =>
                           n13409, C1 => n14683, C2 => n13361, ZN => n12366);
   U12618 : AOI222_X1 port map( A1 => n14698, A2 => n13385, B1 => n14695, B2 =>
                           n13553, C1 => n14692, C2 => n13505, ZN => n12367);
   U12619 : AOI211_X1 port map( C1 => n14719, C2 => n13529, A => n12380, B => 
                           n12381, ZN => n12368);
   U12620 : NAND4_X1 port map( A1 => n12349, A2 => n12350, A3 => n12351, A4 => 
                           n12352, ZN => n1324);
   U12621 : AOI222_X1 port map( A1 => n14689, A2 => n14240, B1 => n14686, B2 =>
                           n13410, C1 => n14683, C2 => n13362, ZN => n12349);
   U12622 : AOI222_X1 port map( A1 => n14698, A2 => n13386, B1 => n14695, B2 =>
                           n13554, C1 => n14692, C2 => n13506, ZN => n12350);
   U12623 : AOI211_X1 port map( C1 => n14719, C2 => n13530, A => n12363, B => 
                           n12364, ZN => n12351);
   U12624 : NAND4_X1 port map( A1 => n12332, A2 => n12333, A3 => n12334, A4 => 
                           n12335, ZN => n1325);
   U12625 : AOI222_X1 port map( A1 => n14689, A2 => n14241, B1 => n14686, B2 =>
                           n13411, C1 => n14683, C2 => n13363, ZN => n12332);
   U12626 : AOI222_X1 port map( A1 => n14698, A2 => n13387, B1 => n14695, B2 =>
                           n13555, C1 => n14692, C2 => n13507, ZN => n12333);
   U12627 : AOI211_X1 port map( C1 => n14719, C2 => n13531, A => n12346, B => 
                           n12347, ZN => n12334);
   U12628 : NAND4_X1 port map( A1 => n12315, A2 => n12316, A3 => n12317, A4 => 
                           n12318, ZN => n1326);
   U12629 : AOI222_X1 port map( A1 => n14689, A2 => n14242, B1 => n14686, B2 =>
                           n13412, C1 => n14683, C2 => n13364, ZN => n12315);
   U12630 : AOI222_X1 port map( A1 => n14698, A2 => n13388, B1 => n14695, B2 =>
                           n13556, C1 => n14692, C2 => n13508, ZN => n12316);
   U12631 : AOI211_X1 port map( C1 => n14719, C2 => n13532, A => n12329, B => 
                           n12330, ZN => n12317);
   U12632 : NAND4_X1 port map( A1 => n12298, A2 => n12299, A3 => n12300, A4 => 
                           n12301, ZN => n1327);
   U12633 : AOI222_X1 port map( A1 => n14689, A2 => n14243, B1 => n14686, B2 =>
                           n13413, C1 => n14683, C2 => n13365, ZN => n12298);
   U12634 : AOI222_X1 port map( A1 => n14698, A2 => n13389, B1 => n14695, B2 =>
                           n13557, C1 => n14692, C2 => n13509, ZN => n12299);
   U12635 : AOI211_X1 port map( C1 => n14719, C2 => n13533, A => n12312, B => 
                           n12313, ZN => n12300);
   U12636 : NAND4_X1 port map( A1 => n12281, A2 => n12282, A3 => n12283, A4 => 
                           n12284, ZN => n1328);
   U12637 : AOI222_X1 port map( A1 => n14689, A2 => n14244, B1 => n14686, B2 =>
                           n13414, C1 => n14683, C2 => n13366, ZN => n12281);
   U12638 : AOI222_X1 port map( A1 => n14698, A2 => n13390, B1 => n14695, B2 =>
                           n13558, C1 => n14692, C2 => n13510, ZN => n12282);
   U12639 : AOI211_X1 port map( C1 => n14719, C2 => n13534, A => n12295, B => 
                           n12296, ZN => n12283);
   U12640 : NAND4_X1 port map( A1 => n12264, A2 => n12265, A3 => n12266, A4 => 
                           n12267, ZN => n1329);
   U12641 : AOI222_X1 port map( A1 => n14689, A2 => n14245, B1 => n14686, B2 =>
                           n13415, C1 => n14683, C2 => n13367, ZN => n12264);
   U12642 : AOI222_X1 port map( A1 => n14698, A2 => n13391, B1 => n14695, B2 =>
                           n13559, C1 => n14692, C2 => n13511, ZN => n12265);
   U12643 : AOI211_X1 port map( C1 => n14719, C2 => n13535, A => n12278, B => 
                           n12279, ZN => n12266);
   U12644 : NAND4_X1 port map( A1 => n12247, A2 => n12248, A3 => n12249, A4 => 
                           n12250, ZN => n1330);
   U12645 : AOI222_X1 port map( A1 => n14689, A2 => n14246, B1 => n14685, B2 =>
                           n13416, C1 => n14682, C2 => n13368, ZN => n12247);
   U12646 : AOI222_X1 port map( A1 => n14698, A2 => n13392, B1 => n14694, B2 =>
                           n13560, C1 => n14691, C2 => n13512, ZN => n12248);
   U12647 : AOI211_X1 port map( C1 => n14719, C2 => n13536, A => n12261, B => 
                           n12262, ZN => n12249);
   U12648 : NAND4_X1 port map( A1 => n12230, A2 => n12231, A3 => n12232, A4 => 
                           n12233, ZN => n1331);
   U12649 : AOI222_X1 port map( A1 => n14689, A2 => n14247, B1 => n14685, B2 =>
                           n13417, C1 => n14682, C2 => n13369, ZN => n12230);
   U12650 : AOI222_X1 port map( A1 => n14698, A2 => n13393, B1 => n14694, B2 =>
                           n13561, C1 => n14691, C2 => n13513, ZN => n12231);
   U12651 : AOI211_X1 port map( C1 => n14719, C2 => n13537, A => n12244, B => 
                           n12245, ZN => n12232);
   U12652 : NAND4_X1 port map( A1 => n12213, A2 => n12214, A3 => n12215, A4 => 
                           n12216, ZN => n1332);
   U12653 : AOI222_X1 port map( A1 => n14689, A2 => n14248, B1 => n14685, B2 =>
                           n13418, C1 => n14682, C2 => n13370, ZN => n12213);
   U12654 : AOI222_X1 port map( A1 => n14698, A2 => n13394, B1 => n14694, B2 =>
                           n13562, C1 => n14691, C2 => n13514, ZN => n12214);
   U12655 : AOI211_X1 port map( C1 => n14719, C2 => n13538, A => n12227, B => 
                           n12228, ZN => n12215);
   U12656 : NAND4_X1 port map( A1 => n12196, A2 => n12197, A3 => n12198, A4 => 
                           n12199, ZN => n1333);
   U12657 : AOI222_X1 port map( A1 => n14689, A2 => n14249, B1 => n14685, B2 =>
                           n13419, C1 => n14682, C2 => n13371, ZN => n12196);
   U12658 : AOI222_X1 port map( A1 => n14698, A2 => n13395, B1 => n14694, B2 =>
                           n13563, C1 => n14691, C2 => n13515, ZN => n12197);
   U12659 : AOI211_X1 port map( C1 => n14719, C2 => n13539, A => n12210, B => 
                           n12211, ZN => n12198);
   U12660 : NAND4_X1 port map( A1 => n12179, A2 => n12180, A3 => n12181, A4 => 
                           n12182, ZN => n1334);
   U12661 : AOI222_X1 port map( A1 => n14690, A2 => n14250, B1 => n14685, B2 =>
                           n13316, C1 => n14682, C2 => n13300, ZN => n12179);
   U12662 : AOI222_X1 port map( A1 => n14699, A2 => n13308, B1 => n14694, B2 =>
                           n13268, C1 => n14691, C2 => n13252, ZN => n12180);
   U12663 : AOI211_X1 port map( C1 => n14720, C2 => n13260, A => n12193, B => 
                           n12194, ZN => n12181);
   U12664 : NAND4_X1 port map( A1 => n12162, A2 => n12163, A3 => n12164, A4 => 
                           n12165, ZN => n1335);
   U12665 : AOI222_X1 port map( A1 => n14690, A2 => n14251, B1 => n14685, B2 =>
                           n13317, C1 => n14682, C2 => n13301, ZN => n12162);
   U12666 : AOI222_X1 port map( A1 => n14699, A2 => n13309, B1 => n14694, B2 =>
                           n13269, C1 => n14691, C2 => n13253, ZN => n12163);
   U12667 : AOI211_X1 port map( C1 => n14720, C2 => n13261, A => n12176, B => 
                           n12177, ZN => n12164);
   U12668 : NAND4_X1 port map( A1 => n12145, A2 => n12146, A3 => n12147, A4 => 
                           n12148, ZN => n1336);
   U12669 : AOI222_X1 port map( A1 => n14690, A2 => n14252, B1 => n14685, B2 =>
                           n13318, C1 => n14682, C2 => n13302, ZN => n12145);
   U12670 : AOI222_X1 port map( A1 => n14699, A2 => n13310, B1 => n14694, B2 =>
                           n13270, C1 => n14691, C2 => n13254, ZN => n12146);
   U12671 : AOI211_X1 port map( C1 => n14720, C2 => n13262, A => n12159, B => 
                           n12160, ZN => n12147);
   U12672 : NAND4_X1 port map( A1 => n12128, A2 => n12129, A3 => n12130, A4 => 
                           n12131, ZN => n1337);
   U12673 : AOI222_X1 port map( A1 => n14690, A2 => n14253, B1 => n14685, B2 =>
                           n13319, C1 => n14682, C2 => n13303, ZN => n12128);
   U12674 : AOI222_X1 port map( A1 => n14699, A2 => n13311, B1 => n14694, B2 =>
                           n13271, C1 => n14691, C2 => n13255, ZN => n12129);
   U12675 : AOI211_X1 port map( C1 => n14720, C2 => n13263, A => n12142, B => 
                           n12143, ZN => n12130);
   U12676 : NAND4_X1 port map( A1 => n12111, A2 => n12112, A3 => n12113, A4 => 
                           n12114, ZN => n1338);
   U12677 : AOI222_X1 port map( A1 => n14690, A2 => n14254, B1 => n14685, B2 =>
                           n13320, C1 => n14682, C2 => n13304, ZN => n12111);
   U12678 : AOI222_X1 port map( A1 => n14699, A2 => n13312, B1 => n14694, B2 =>
                           n13272, C1 => n14691, C2 => n13256, ZN => n12112);
   U12679 : AOI211_X1 port map( C1 => n14720, C2 => n13264, A => n12125, B => 
                           n12126, ZN => n12113);
   U12680 : NAND4_X1 port map( A1 => n12094, A2 => n12095, A3 => n12096, A4 => 
                           n12097, ZN => n1339);
   U12681 : AOI222_X1 port map( A1 => n14690, A2 => n14255, B1 => n14685, B2 =>
                           n13321, C1 => n14682, C2 => n13305, ZN => n12094);
   U12682 : AOI222_X1 port map( A1 => n14699, A2 => n13313, B1 => n14694, B2 =>
                           n13273, C1 => n14691, C2 => n13257, ZN => n12095);
   U12683 : AOI211_X1 port map( C1 => n14720, C2 => n13265, A => n12108, B => 
                           n12109, ZN => n12096);
   U12684 : NAND4_X1 port map( A1 => n12077, A2 => n12078, A3 => n12079, A4 => 
                           n12080, ZN => n1340);
   U12685 : AOI222_X1 port map( A1 => n14690, A2 => n14256, B1 => n14685, B2 =>
                           n13322, C1 => n14682, C2 => n13306, ZN => n12077);
   U12686 : AOI222_X1 port map( A1 => n14699, A2 => n13314, B1 => n14694, B2 =>
                           n13274, C1 => n14691, C2 => n13258, ZN => n12078);
   U12687 : AOI211_X1 port map( C1 => n14720, C2 => n13266, A => n12091, B => 
                           n12092, ZN => n12079);
   U12688 : NAND4_X1 port map( A1 => n12026, A2 => n12027, A3 => n12028, A4 => 
                           n12029, ZN => n1341);
   U12689 : AOI222_X1 port map( A1 => n14690, A2 => n14257, B1 => n14685, B2 =>
                           n13323, C1 => n14682, C2 => n13307, ZN => n12026);
   U12690 : AOI222_X1 port map( A1 => n14699, A2 => n13315, B1 => n14694, B2 =>
                           n13275, C1 => n14691, C2 => n13259, ZN => n12027);
   U12691 : AOI211_X1 port map( C1 => n14720, C2 => n13267, A => n12062, B => 
                           n12063, ZN => n12028);
   U12692 : OAI22_X1 port map( A1 => n14954, A2 => n15062, B1 => n14953, B2 => 
                           n14482, ZN => n1950);
   U12693 : OAI22_X1 port map( A1 => n14954, A2 => n15065, B1 => n14953, B2 => 
                           n14483, ZN => n1951);
   U12694 : OAI22_X1 port map( A1 => n14954, A2 => n15068, B1 => n14953, B2 => 
                           n14484, ZN => n1952);
   U12695 : OAI22_X1 port map( A1 => n14954, A2 => n15071, B1 => n14953, B2 => 
                           n14485, ZN => n1953);
   U12696 : OAI22_X1 port map( A1 => n14954, A2 => n15074, B1 => n14953, B2 => 
                           n14486, ZN => n1954);
   U12697 : OAI22_X1 port map( A1 => n14955, A2 => n15077, B1 => n14953, B2 => 
                           n14487, ZN => n1955);
   U12698 : OAI22_X1 port map( A1 => n14955, A2 => n15080, B1 => n14953, B2 => 
                           n14488, ZN => n1956);
   U12699 : OAI22_X1 port map( A1 => n14955, A2 => n15083, B1 => n14953, B2 => 
                           n14489, ZN => n1957);
   U12700 : OAI22_X1 port map( A1 => n14955, A2 => n15086, B1 => n14953, B2 => 
                           n14490, ZN => n1958);
   U12701 : OAI22_X1 port map( A1 => n14955, A2 => n15089, B1 => n14953, B2 => 
                           n14491, ZN => n1959);
   U12702 : OAI22_X1 port map( A1 => n14956, A2 => n15092, B1 => n14953, B2 => 
                           n14492, ZN => n1960);
   U12703 : OAI22_X1 port map( A1 => n14956, A2 => n15095, B1 => n14953, B2 => 
                           n14493, ZN => n1961);
   U12704 : OAI22_X1 port map( A1 => n14956, A2 => n15098, B1 => n12000, B2 => 
                           n14494, ZN => n1962);
   U12705 : OAI22_X1 port map( A1 => n14956, A2 => n15101, B1 => n12000, B2 => 
                           n14495, ZN => n1963);
   U12706 : OAI22_X1 port map( A1 => n14956, A2 => n15104, B1 => n12000, B2 => 
                           n14496, ZN => n1964);
   U12707 : OAI22_X1 port map( A1 => n14957, A2 => n15107, B1 => n14953, B2 => 
                           n14497, ZN => n1965);
   U12708 : OAI22_X1 port map( A1 => n14957, A2 => n15110, B1 => n14953, B2 => 
                           n14498, ZN => n1966);
   U12709 : OAI22_X1 port map( A1 => n14957, A2 => n15113, B1 => n14953, B2 => 
                           n14499, ZN => n1967);
   U12710 : OAI22_X1 port map( A1 => n14957, A2 => n15116, B1 => n14953, B2 => 
                           n14500, ZN => n1968);
   U12711 : OAI22_X1 port map( A1 => n14957, A2 => n15119, B1 => n14953, B2 => 
                           n14501, ZN => n1969);
   U12712 : OAI22_X1 port map( A1 => n14958, A2 => n15122, B1 => n14953, B2 => 
                           n14502, ZN => n1970);
   U12713 : OAI22_X1 port map( A1 => n14958, A2 => n15125, B1 => n14953, B2 => 
                           n14503, ZN => n1971);
   U12714 : OAI22_X1 port map( A1 => n14958, A2 => n15128, B1 => n14953, B2 => 
                           n14504, ZN => n1972);
   U12715 : OAI22_X1 port map( A1 => n14958, A2 => n15131, B1 => n14953, B2 => 
                           n14505, ZN => n1973);
   U12716 : OAI22_X1 port map( A1 => n15026, A2 => n15061, B1 => n15025, B2 => 
                           n14506, ZN => n2206);
   U12717 : OAI22_X1 port map( A1 => n15026, A2 => n15064, B1 => n15025, B2 => 
                           n14507, ZN => n2207);
   U12718 : OAI22_X1 port map( A1 => n15026, A2 => n15067, B1 => n15025, B2 => 
                           n14508, ZN => n2208);
   U12719 : OAI22_X1 port map( A1 => n15026, A2 => n15070, B1 => n15025, B2 => 
                           n14509, ZN => n2209);
   U12720 : OAI22_X1 port map( A1 => n15026, A2 => n15073, B1 => n15025, B2 => 
                           n14510, ZN => n2210);
   U12721 : OAI22_X1 port map( A1 => n15027, A2 => n15076, B1 => n15025, B2 => 
                           n14511, ZN => n2211);
   U12722 : OAI22_X1 port map( A1 => n15027, A2 => n15079, B1 => n15025, B2 => 
                           n14512, ZN => n2212);
   U12723 : OAI22_X1 port map( A1 => n15027, A2 => n15082, B1 => n15025, B2 => 
                           n14513, ZN => n2213);
   U12724 : OAI22_X1 port map( A1 => n15027, A2 => n15085, B1 => n15025, B2 => 
                           n14514, ZN => n2214);
   U12725 : OAI22_X1 port map( A1 => n15027, A2 => n15088, B1 => n15025, B2 => 
                           n14515, ZN => n2215);
   U12726 : OAI22_X1 port map( A1 => n15028, A2 => n15091, B1 => n15025, B2 => 
                           n14516, ZN => n2216);
   U12727 : OAI22_X1 port map( A1 => n15028, A2 => n15094, B1 => n15025, B2 => 
                           n14517, ZN => n2217);
   U12728 : OAI22_X1 port map( A1 => n15028, A2 => n15097, B1 => n11990, B2 => 
                           n14518, ZN => n2218);
   U12729 : OAI22_X1 port map( A1 => n15028, A2 => n15100, B1 => n11990, B2 => 
                           n14519, ZN => n2219);
   U12730 : OAI22_X1 port map( A1 => n15028, A2 => n15103, B1 => n11990, B2 => 
                           n14520, ZN => n2220);
   U12731 : OAI22_X1 port map( A1 => n15029, A2 => n15106, B1 => n15025, B2 => 
                           n14521, ZN => n2221);
   U12732 : OAI22_X1 port map( A1 => n15029, A2 => n15109, B1 => n15025, B2 => 
                           n14522, ZN => n2222);
   U12733 : OAI22_X1 port map( A1 => n15029, A2 => n15112, B1 => n15025, B2 => 
                           n14523, ZN => n2223);
   U12734 : OAI22_X1 port map( A1 => n15029, A2 => n15115, B1 => n15025, B2 => 
                           n14524, ZN => n2224);
   U12735 : OAI22_X1 port map( A1 => n15029, A2 => n15118, B1 => n15025, B2 => 
                           n14525, ZN => n2225);
   U12736 : OAI22_X1 port map( A1 => n15030, A2 => n15121, B1 => n15025, B2 => 
                           n14526, ZN => n2226);
   U12737 : OAI22_X1 port map( A1 => n15030, A2 => n15124, B1 => n15025, B2 => 
                           n14527, ZN => n2227);
   U12738 : OAI22_X1 port map( A1 => n15030, A2 => n15127, B1 => n15025, B2 => 
                           n14528, ZN => n2228);
   U12739 : OAI22_X1 port map( A1 => n15030, A2 => n15130, B1 => n15025, B2 => 
                           n14529, ZN => n2229);
   U12740 : NAND2_X1 port map( A1 => ADD_WR(1), A2 => ADD_WR(0), ZN => n11988);
   U12741 : NAND2_X1 port map( A1 => ADD_WR(1), A2 => n10991, ZN => n11986);
   U12742 : NAND2_X1 port map( A1 => ADD_WR(0), A2 => n10990, ZN => n11984);
   U12743 : NOR3_X1 port map( A1 => ADD_RD2(2), A2 => ADD_RD2(4), A3 => n11004,
                           ZN => n12624);
   U12744 : NOR3_X1 port map( A1 => n11005, A2 => ADD_RD2(4), A3 => n11004, ZN 
                           => n12629);
   U12745 : NOR3_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), A3 => n11005,
                           ZN => n12630);
   U12746 : NOR3_X1 port map( A1 => ADD_RD1(2), A2 => ADD_RD1(4), A3 => n10996,
                           ZN => n12043);
   U12747 : NOR3_X1 port map( A1 => n10997, A2 => ADD_RD1(4), A3 => n10996, ZN 
                           => n12048);
   U12748 : NOR3_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), A3 => n10997,
                           ZN => n12049);
   U12749 : NOR3_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), A3 => 
                           ADD_RD2(2), ZN => n12625);
   U12750 : NOR3_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), A3 => 
                           ADD_RD1(2), ZN => n12044);
   U12751 : AND3_X1 port map( A1 => n14678, A2 => n11007, A3 => ADD_RD2(1), ZN 
                           => n13181);
   U12752 : AND3_X1 port map( A1 => n14776, A2 => n10999, A3 => ADD_RD1(1), ZN 
                           => n12600);
   U12753 : AND3_X1 port map( A1 => n14678, A2 => n11006, A3 => ADD_RD2(0), ZN 
                           => n13183);
   U12754 : AND3_X1 port map( A1 => n14776, A2 => n10998, A3 => ADD_RD1(0), ZN 
                           => n12602);
   U12755 : INV_X1 port map( A => RESET, ZN => n10986);
   U12756 : AND2_X1 port map( A1 => RD2, A2 => ENABLE, ZN => n12616);
   U12757 : AND2_X1 port map( A1 => RD1, A2 => ENABLE, ZN => n12035);
   U12758 : AND3_X1 port map( A1 => ADD_RD2(0), A2 => n14678, A3 => ADD_RD2(1),
                           ZN => n12620);
   U12759 : AND3_X1 port map( A1 => ADD_RD1(0), A2 => n14776, A3 => ADD_RD1(1),
                           ZN => n12039);
   U12760 : NAND2_X1 port map( A1 => DATAIN(8), A2 => n15167, ZN => n11972);
   U12761 : NAND2_X1 port map( A1 => DATAIN(9), A2 => n15167, ZN => n11971);
   U12762 : NAND2_X1 port map( A1 => DATAIN(10), A2 => n15167, ZN => n11970);
   U12763 : NAND2_X1 port map( A1 => DATAIN(11), A2 => n15167, ZN => n11969);
   U12764 : NAND2_X1 port map( A1 => DATAIN(12), A2 => n15167, ZN => n11968);
   U12765 : NAND2_X1 port map( A1 => DATAIN(13), A2 => n15167, ZN => n11967);
   U12766 : NAND2_X1 port map( A1 => DATAIN(14), A2 => n15167, ZN => n11966);
   U12767 : NAND2_X1 port map( A1 => DATAIN(15), A2 => n15167, ZN => n11965);
   U12768 : NAND2_X1 port map( A1 => DATAIN(16), A2 => n15167, ZN => n11964);
   U12769 : NAND2_X1 port map( A1 => DATAIN(17), A2 => n15167, ZN => n11963);
   U12770 : NAND2_X1 port map( A1 => DATAIN(18), A2 => n15167, ZN => n11962);
   U12771 : NAND2_X1 port map( A1 => DATAIN(19), A2 => n15167, ZN => n11961);
   U12772 : NAND2_X1 port map( A1 => DATAIN(20), A2 => n15166, ZN => n11960);
   U12773 : NAND2_X1 port map( A1 => DATAIN(21), A2 => n15166, ZN => n11959);
   U12774 : NAND2_X1 port map( A1 => DATAIN(22), A2 => n15166, ZN => n11958);
   U12775 : NAND2_X1 port map( A1 => DATAIN(23), A2 => n15166, ZN => n11957);
   U12776 : NAND2_X1 port map( A1 => DATAIN(24), A2 => n15166, ZN => n11956);
   U12777 : NAND2_X1 port map( A1 => DATAIN(25), A2 => n15166, ZN => n11955);
   U12778 : NAND2_X1 port map( A1 => DATAIN(26), A2 => n15166, ZN => n11954);
   U12779 : NAND2_X1 port map( A1 => DATAIN(27), A2 => n15166, ZN => n11953);
   U12780 : NAND2_X1 port map( A1 => DATAIN(28), A2 => n15166, ZN => n11952);
   U12781 : NAND2_X1 port map( A1 => DATAIN(29), A2 => n15166, ZN => n11951);
   U12782 : NAND2_X1 port map( A1 => DATAIN(30), A2 => n15166, ZN => n11950);
   U12783 : NAND2_X1 port map( A1 => DATAIN(31), A2 => n15166, ZN => n11948);
   U12784 : NAND2_X1 port map( A1 => DATAIN(0), A2 => n15168, ZN => n11980);
   U12785 : NAND2_X1 port map( A1 => DATAIN(1), A2 => n15168, ZN => n11979);
   U12786 : NAND2_X1 port map( A1 => DATAIN(2), A2 => n15168, ZN => n11978);
   U12787 : NAND2_X1 port map( A1 => DATAIN(3), A2 => n15168, ZN => n11977);
   U12788 : NAND2_X1 port map( A1 => DATAIN(4), A2 => n15168, ZN => n11976);
   U12789 : NAND2_X1 port map( A1 => DATAIN(5), A2 => n15168, ZN => n11975);
   U12790 : NAND2_X1 port map( A1 => DATAIN(6), A2 => n15168, ZN => n11974);
   U12791 : NAND2_X1 port map( A1 => DATAIN(7), A2 => n15168, ZN => n11973);
   U12792 : INV_X1 port map( A => ADD_RD2(3), ZN => n11004);
   U12793 : INV_X1 port map( A => ADD_RD1(3), ZN => n10996);
   U12794 : INV_X1 port map( A => ADD_RD2(2), ZN => n11005);
   U12795 : INV_X1 port map( A => ADD_RD1(2), ZN => n10997);
   U12796 : AND3_X1 port map( A1 => n11005, A2 => n11004, A3 => ADD_RD2(4), ZN 
                           => n14578);
   U12797 : AND3_X1 port map( A1 => n10997, A2 => n10996, A3 => ADD_RD1(4), ZN 
                           => n14579);
   U12798 : AND3_X1 port map( A1 => ADD_RD2(2), A2 => n11004, A3 => ADD_RD2(4),
                           ZN => n14580);
   U12799 : AND3_X1 port map( A1 => ADD_RD1(2), A2 => n10996, A3 => ADD_RD1(4),
                           ZN => n14581);
   U12800 : AND3_X1 port map( A1 => WR, A2 => ENABLE, A3 => ADD_WR(4), ZN => 
                           n12010);
   U12801 : AND3_X1 port map( A1 => ENABLE, A2 => n10987, A3 => WR, ZN => 
                           n11989);
   U12802 : INV_X1 port map( A => ADD_WR(4), ZN => n10987);
   U12803 : AND3_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(2), A3 => 
                           ADD_RD2(4), ZN => n14582);
   U12804 : AND3_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(2), A3 => 
                           ADD_RD1(4), ZN => n14583);
   U12805 : INV_X1 port map( A => ADD_WR(3), ZN => n10988);
   U12806 : INV_X1 port map( A => ADD_WR(2), ZN => n10989);
   U12807 : INV_X1 port map( A => ADD_WR(0), ZN => n10991);
   U12808 : INV_X1 port map( A => ADD_WR(1), ZN => n10990);
   U12809 : INV_X1 port map( A => ADD_RD2(1), ZN => n11006);
   U12810 : INV_X1 port map( A => ADD_RD1(1), ZN => n10998);
   U12811 : INV_X1 port map( A => ADD_RD2(0), ZN => n11007);
   U12812 : INV_X1 port map( A => ADD_RD1(0), ZN => n10999);
   U12813 : INV_X1 port map( A => n14582, ZN => n14662);
   U12814 : INV_X1 port map( A => n14583, ZN => n14760);
   U12815 : CLKBUF_X1 port map( A => n10986, Z => n15171);

end SYN_Beh;
