
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_BOOTHMUL_NBIT8 is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_BOOTHMUL_NBIT8;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity SETTLER_NBIT16_0_DW01_inc_0 is

   port( A : in std_logic_vector (15 downto 0);  SUM : out std_logic_vector (15
         downto 0));

end SETTLER_NBIT16_0_DW01_inc_0;

architecture SYN_rpl of SETTLER_NBIT16_0_DW01_inc_0 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component HA_X1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_15_port, carry_14_port, carry_13_port, carry_12_port, 
      carry_11_port, carry_10_port, carry_9_port, carry_8_port, carry_7_port, 
      carry_6_port, carry_5_port, carry_4_port, carry_3_port : std_logic;

begin
   
   U1_1_14 : HA_X1 port map( A => A(14), B => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_1_13 : HA_X1 port map( A => A(13), B => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_1_12 : HA_X1 port map( A => A(12), B => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_1_11 : HA_X1 port map( A => A(11), B => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_1_10 : HA_X1 port map( A => A(10), B => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_1_9 : HA_X1 port map( A => A(9), B => carry_9_port, CO => carry_10_port, 
                           S => SUM(9));
   U1_1_8 : HA_X1 port map( A => A(8), B => carry_8_port, CO => carry_9_port, S
                           => SUM(8));
   U1_1_7 : HA_X1 port map( A => A(7), B => carry_7_port, CO => carry_8_port, S
                           => SUM(7));
   U1_1_6 : HA_X1 port map( A => A(6), B => carry_6_port, CO => carry_7_port, S
                           => SUM(6));
   U1_1_5 : HA_X1 port map( A => A(5), B => carry_5_port, CO => carry_6_port, S
                           => SUM(5));
   U1_1_4 : HA_X1 port map( A => A(4), B => carry_4_port, CO => carry_5_port, S
                           => SUM(4));
   U1_1_3 : HA_X1 port map( A => A(3), B => carry_3_port, CO => carry_4_port, S
                           => SUM(3));
   U1_1_2 : HA_X1 port map( A => A(2), B => A(1), CO => carry_3_port, S => 
                           SUM(2));
   U1 : INV_X1 port map( A => A(1), ZN => SUM(1));
   U2 : XOR2_X1 port map( A => carry_15_port, B => A(15), Z => SUM(15));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity SETTLER_NBIT16_3_DW01_inc_0 is

   port( A : in std_logic_vector (15 downto 0);  SUM : out std_logic_vector (15
         downto 0));

end SETTLER_NBIT16_3_DW01_inc_0;

architecture SYN_rpl of SETTLER_NBIT16_3_DW01_inc_0 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component HA_X1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_15_port, carry_14_port, carry_13_port, carry_12_port, 
      carry_11_port, carry_10_port, carry_9_port, carry_8_port, carry_7_port, 
      carry_6_port, carry_5_port, carry_4_port, carry_3_port : std_logic;

begin
   
   U1_1_14 : HA_X1 port map( A => A(14), B => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_1_13 : HA_X1 port map( A => A(13), B => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_1_12 : HA_X1 port map( A => A(12), B => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_1_11 : HA_X1 port map( A => A(11), B => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_1_10 : HA_X1 port map( A => A(10), B => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_1_9 : HA_X1 port map( A => A(9), B => carry_9_port, CO => carry_10_port, 
                           S => SUM(9));
   U1_1_8 : HA_X1 port map( A => A(8), B => carry_8_port, CO => carry_9_port, S
                           => SUM(8));
   U1_1_7 : HA_X1 port map( A => A(7), B => carry_7_port, CO => carry_8_port, S
                           => SUM(7));
   U1_1_6 : HA_X1 port map( A => A(6), B => carry_6_port, CO => carry_7_port, S
                           => SUM(6));
   U1_1_5 : HA_X1 port map( A => A(5), B => carry_5_port, CO => carry_6_port, S
                           => SUM(5));
   U1_1_4 : HA_X1 port map( A => A(4), B => carry_4_port, CO => carry_5_port, S
                           => SUM(4));
   U1_1_3 : HA_X1 port map( A => A(3), B => carry_3_port, CO => carry_4_port, S
                           => SUM(3));
   U1_1_2 : HA_X1 port map( A => A(2), B => A(1), CO => carry_3_port, S => 
                           SUM(2));
   U1 : INV_X1 port map( A => A(1), ZN => SUM(1));
   U2 : XOR2_X1 port map( A => carry_15_port, B => A(15), Z => SUM(15));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity SETTLER_NBIT16_2_DW01_inc_0 is

   port( A : in std_logic_vector (15 downto 0);  SUM : out std_logic_vector (15
         downto 0));

end SETTLER_NBIT16_2_DW01_inc_0;

architecture SYN_rpl of SETTLER_NBIT16_2_DW01_inc_0 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component HA_X1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_15_port, carry_14_port, carry_13_port, carry_12_port, 
      carry_11_port, carry_10_port, carry_9_port, carry_8_port, carry_7_port, 
      carry_6_port, carry_5_port, carry_4_port, carry_3_port : std_logic;

begin
   
   U1_1_14 : HA_X1 port map( A => A(14), B => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_1_13 : HA_X1 port map( A => A(13), B => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_1_12 : HA_X1 port map( A => A(12), B => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_1_11 : HA_X1 port map( A => A(11), B => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_1_10 : HA_X1 port map( A => A(10), B => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_1_9 : HA_X1 port map( A => A(9), B => carry_9_port, CO => carry_10_port, 
                           S => SUM(9));
   U1_1_8 : HA_X1 port map( A => A(8), B => carry_8_port, CO => carry_9_port, S
                           => SUM(8));
   U1_1_7 : HA_X1 port map( A => A(7), B => carry_7_port, CO => carry_8_port, S
                           => SUM(7));
   U1_1_6 : HA_X1 port map( A => A(6), B => carry_6_port, CO => carry_7_port, S
                           => SUM(6));
   U1_1_5 : HA_X1 port map( A => A(5), B => carry_5_port, CO => carry_6_port, S
                           => SUM(5));
   U1_1_4 : HA_X1 port map( A => A(4), B => carry_4_port, CO => carry_5_port, S
                           => SUM(4));
   U1_1_3 : HA_X1 port map( A => A(3), B => carry_3_port, CO => carry_4_port, S
                           => SUM(3));
   U1_1_2 : HA_X1 port map( A => A(2), B => A(1), CO => carry_3_port, S => 
                           SUM(2));
   U1 : INV_X1 port map( A => A(1), ZN => SUM(1));
   U2 : XOR2_X1 port map( A => carry_15_port, B => A(15), Z => SUM(15));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity SETTLER_NBIT16_1_DW01_inc_0 is

   port( A : in std_logic_vector (15 downto 0);  SUM : out std_logic_vector (15
         downto 0));

end SETTLER_NBIT16_1_DW01_inc_0;

architecture SYN_rpl of SETTLER_NBIT16_1_DW01_inc_0 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component HA_X1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_15_port, carry_14_port, carry_13_port, carry_12_port, 
      carry_11_port, carry_10_port, carry_9_port, carry_8_port, carry_7_port, 
      carry_6_port, carry_5_port, carry_4_port, carry_3_port : std_logic;

begin
   
   U1_1_14 : HA_X1 port map( A => A(14), B => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_1_13 : HA_X1 port map( A => A(13), B => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_1_12 : HA_X1 port map( A => A(12), B => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_1_11 : HA_X1 port map( A => A(11), B => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_1_10 : HA_X1 port map( A => A(10), B => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_1_9 : HA_X1 port map( A => A(9), B => carry_9_port, CO => carry_10_port, 
                           S => SUM(9));
   U1_1_8 : HA_X1 port map( A => A(8), B => carry_8_port, CO => carry_9_port, S
                           => SUM(8));
   U1_1_7 : HA_X1 port map( A => A(7), B => carry_7_port, CO => carry_8_port, S
                           => SUM(7));
   U1_1_6 : HA_X1 port map( A => A(6), B => carry_6_port, CO => carry_7_port, S
                           => SUM(6));
   U1_1_5 : HA_X1 port map( A => A(5), B => carry_5_port, CO => carry_6_port, S
                           => SUM(5));
   U1_1_4 : HA_X1 port map( A => A(4), B => carry_4_port, CO => carry_5_port, S
                           => SUM(4));
   U1_1_3 : HA_X1 port map( A => A(3), B => carry_3_port, CO => carry_4_port, S
                           => SUM(3));
   U1_1_2 : HA_X1 port map( A => A(2), B => A(1), CO => carry_3_port, S => 
                           SUM(2));
   U1 : INV_X1 port map( A => A(1), ZN => SUM(1));
   U2 : XOR2_X1 port map( A => carry_15_port, B => A(15), Z => SUM(15));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_767 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_767;

architecture SYN_ARCH2 of ND2_767 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_766 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_766;

architecture SYN_ARCH2 of ND2_766 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_765 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_765;

architecture SYN_ARCH2 of ND2_765 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_764 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_764;

architecture SYN_ARCH2 of ND2_764 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_763 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_763;

architecture SYN_ARCH2 of ND2_763 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_762 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_762;

architecture SYN_ARCH2 of ND2_762 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_761 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_761;

architecture SYN_ARCH2 of ND2_761 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_760 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_760;

architecture SYN_ARCH2 of ND2_760 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_759 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_759;

architecture SYN_ARCH2 of ND2_759 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_758 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_758;

architecture SYN_ARCH2 of ND2_758 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_757 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_757;

architecture SYN_ARCH2 of ND2_757 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_756 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_756;

architecture SYN_ARCH2 of ND2_756 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_755 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_755;

architecture SYN_ARCH2 of ND2_755 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_754 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_754;

architecture SYN_ARCH2 of ND2_754 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_753 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_753;

architecture SYN_ARCH2 of ND2_753 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_752 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_752;

architecture SYN_ARCH2 of ND2_752 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_751 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_751;

architecture SYN_ARCH2 of ND2_751 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_750 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_750;

architecture SYN_ARCH2 of ND2_750 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_749 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_749;

architecture SYN_ARCH2 of ND2_749 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_748 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_748;

architecture SYN_ARCH2 of ND2_748 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_747 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_747;

architecture SYN_ARCH2 of ND2_747 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_746 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_746;

architecture SYN_ARCH2 of ND2_746 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_745 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_745;

architecture SYN_ARCH2 of ND2_745 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_744 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_744;

architecture SYN_ARCH2 of ND2_744 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_743 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_743;

architecture SYN_ARCH2 of ND2_743 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_742 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_742;

architecture SYN_ARCH2 of ND2_742 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_741 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_741;

architecture SYN_ARCH2 of ND2_741 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_740 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_740;

architecture SYN_ARCH2 of ND2_740 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_739 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_739;

architecture SYN_ARCH2 of ND2_739 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_738 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_738;

architecture SYN_ARCH2 of ND2_738 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_737 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_737;

architecture SYN_ARCH2 of ND2_737 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_736 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_736;

architecture SYN_ARCH2 of ND2_736 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_735 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_735;

architecture SYN_ARCH2 of ND2_735 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_734 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_734;

architecture SYN_ARCH2 of ND2_734 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_733 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_733;

architecture SYN_ARCH2 of ND2_733 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_732 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_732;

architecture SYN_ARCH2 of ND2_732 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_731 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_731;

architecture SYN_ARCH2 of ND2_731 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_730 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_730;

architecture SYN_ARCH2 of ND2_730 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_729 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_729;

architecture SYN_ARCH2 of ND2_729 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_728 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_728;

architecture SYN_ARCH2 of ND2_728 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_727 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_727;

architecture SYN_ARCH2 of ND2_727 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_726 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_726;

architecture SYN_ARCH2 of ND2_726 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_725 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_725;

architecture SYN_ARCH2 of ND2_725 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_724 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_724;

architecture SYN_ARCH2 of ND2_724 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_723 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_723;

architecture SYN_ARCH2 of ND2_723 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_722 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_722;

architecture SYN_ARCH2 of ND2_722 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_721 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_721;

architecture SYN_ARCH2 of ND2_721 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_720 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_720;

architecture SYN_ARCH2 of ND2_720 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_719 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_719;

architecture SYN_ARCH2 of ND2_719 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_718 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_718;

architecture SYN_ARCH2 of ND2_718 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_717 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_717;

architecture SYN_ARCH2 of ND2_717 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_716 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_716;

architecture SYN_ARCH2 of ND2_716 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_715 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_715;

architecture SYN_ARCH2 of ND2_715 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_714 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_714;

architecture SYN_ARCH2 of ND2_714 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_713 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_713;

architecture SYN_ARCH2 of ND2_713 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_712 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_712;

architecture SYN_ARCH2 of ND2_712 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_711 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_711;

architecture SYN_ARCH2 of ND2_711 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_710 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_710;

architecture SYN_ARCH2 of ND2_710 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_709 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_709;

architecture SYN_ARCH2 of ND2_709 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_708 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_708;

architecture SYN_ARCH2 of ND2_708 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_707 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_707;

architecture SYN_ARCH2 of ND2_707 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_706 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_706;

architecture SYN_ARCH2 of ND2_706 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_705 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_705;

architecture SYN_ARCH2 of ND2_705 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_704 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_704;

architecture SYN_ARCH2 of ND2_704 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_703 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_703;

architecture SYN_ARCH2 of ND2_703 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_702 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_702;

architecture SYN_ARCH2 of ND2_702 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_701 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_701;

architecture SYN_ARCH2 of ND2_701 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_700 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_700;

architecture SYN_ARCH2 of ND2_700 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_699 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_699;

architecture SYN_ARCH2 of ND2_699 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_698 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_698;

architecture SYN_ARCH2 of ND2_698 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_697 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_697;

architecture SYN_ARCH2 of ND2_697 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_696 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_696;

architecture SYN_ARCH2 of ND2_696 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_695 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_695;

architecture SYN_ARCH2 of ND2_695 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_694 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_694;

architecture SYN_ARCH2 of ND2_694 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_693 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_693;

architecture SYN_ARCH2 of ND2_693 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_692 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_692;

architecture SYN_ARCH2 of ND2_692 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_691 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_691;

architecture SYN_ARCH2 of ND2_691 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_690 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_690;

architecture SYN_ARCH2 of ND2_690 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_689 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_689;

architecture SYN_ARCH2 of ND2_689 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_688 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_688;

architecture SYN_ARCH2 of ND2_688 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_687 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_687;

architecture SYN_ARCH2 of ND2_687 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_686 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_686;

architecture SYN_ARCH2 of ND2_686 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_685 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_685;

architecture SYN_ARCH2 of ND2_685 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_684 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_684;

architecture SYN_ARCH2 of ND2_684 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_683 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_683;

architecture SYN_ARCH2 of ND2_683 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_682 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_682;

architecture SYN_ARCH2 of ND2_682 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_681 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_681;

architecture SYN_ARCH2 of ND2_681 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_680 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_680;

architecture SYN_ARCH2 of ND2_680 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_679 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_679;

architecture SYN_ARCH2 of ND2_679 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_678 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_678;

architecture SYN_ARCH2 of ND2_678 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_677 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_677;

architecture SYN_ARCH2 of ND2_677 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_676 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_676;

architecture SYN_ARCH2 of ND2_676 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_675 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_675;

architecture SYN_ARCH2 of ND2_675 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_674 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_674;

architecture SYN_ARCH2 of ND2_674 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_673 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_673;

architecture SYN_ARCH2 of ND2_673 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_672 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_672;

architecture SYN_ARCH2 of ND2_672 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_671 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_671;

architecture SYN_ARCH2 of ND2_671 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_670 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_670;

architecture SYN_ARCH2 of ND2_670 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_669 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_669;

architecture SYN_ARCH2 of ND2_669 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_668 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_668;

architecture SYN_ARCH2 of ND2_668 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_667 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_667;

architecture SYN_ARCH2 of ND2_667 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_666 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_666;

architecture SYN_ARCH2 of ND2_666 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_665 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_665;

architecture SYN_ARCH2 of ND2_665 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_664 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_664;

architecture SYN_ARCH2 of ND2_664 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_663 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_663;

architecture SYN_ARCH2 of ND2_663 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_662 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_662;

architecture SYN_ARCH2 of ND2_662 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_661 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_661;

architecture SYN_ARCH2 of ND2_661 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_660 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_660;

architecture SYN_ARCH2 of ND2_660 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_659 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_659;

architecture SYN_ARCH2 of ND2_659 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_658 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_658;

architecture SYN_ARCH2 of ND2_658 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_657 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_657;

architecture SYN_ARCH2 of ND2_657 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_656 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_656;

architecture SYN_ARCH2 of ND2_656 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_655 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_655;

architecture SYN_ARCH2 of ND2_655 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_654 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_654;

architecture SYN_ARCH2 of ND2_654 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_653 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_653;

architecture SYN_ARCH2 of ND2_653 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_652 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_652;

architecture SYN_ARCH2 of ND2_652 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_651 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_651;

architecture SYN_ARCH2 of ND2_651 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_650 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_650;

architecture SYN_ARCH2 of ND2_650 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_649 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_649;

architecture SYN_ARCH2 of ND2_649 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_648 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_648;

architecture SYN_ARCH2 of ND2_648 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_647 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_647;

architecture SYN_ARCH2 of ND2_647 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_646 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_646;

architecture SYN_ARCH2 of ND2_646 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_645 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_645;

architecture SYN_ARCH2 of ND2_645 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_644 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_644;

architecture SYN_ARCH2 of ND2_644 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_643 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_643;

architecture SYN_ARCH2 of ND2_643 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_642 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_642;

architecture SYN_ARCH2 of ND2_642 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_641 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_641;

architecture SYN_ARCH2 of ND2_641 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_640 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_640;

architecture SYN_ARCH2 of ND2_640 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_639 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_639;

architecture SYN_ARCH2 of ND2_639 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_638 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_638;

architecture SYN_ARCH2 of ND2_638 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_637 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_637;

architecture SYN_ARCH2 of ND2_637 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_636 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_636;

architecture SYN_ARCH2 of ND2_636 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_635 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_635;

architecture SYN_ARCH2 of ND2_635 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_634 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_634;

architecture SYN_ARCH2 of ND2_634 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_633 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_633;

architecture SYN_ARCH2 of ND2_633 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_632 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_632;

architecture SYN_ARCH2 of ND2_632 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_631 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_631;

architecture SYN_ARCH2 of ND2_631 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_630 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_630;

architecture SYN_ARCH2 of ND2_630 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_629 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_629;

architecture SYN_ARCH2 of ND2_629 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_628 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_628;

architecture SYN_ARCH2 of ND2_628 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_627 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_627;

architecture SYN_ARCH2 of ND2_627 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_626 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_626;

architecture SYN_ARCH2 of ND2_626 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_625 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_625;

architecture SYN_ARCH2 of ND2_625 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_624 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_624;

architecture SYN_ARCH2 of ND2_624 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_623 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_623;

architecture SYN_ARCH2 of ND2_623 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_622 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_622;

architecture SYN_ARCH2 of ND2_622 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_621 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_621;

architecture SYN_ARCH2 of ND2_621 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_620 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_620;

architecture SYN_ARCH2 of ND2_620 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_619 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_619;

architecture SYN_ARCH2 of ND2_619 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_618 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_618;

architecture SYN_ARCH2 of ND2_618 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_617 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_617;

architecture SYN_ARCH2 of ND2_617 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_616 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_616;

architecture SYN_ARCH2 of ND2_616 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_615 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_615;

architecture SYN_ARCH2 of ND2_615 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_614 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_614;

architecture SYN_ARCH2 of ND2_614 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_613 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_613;

architecture SYN_ARCH2 of ND2_613 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_612 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_612;

architecture SYN_ARCH2 of ND2_612 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_611 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_611;

architecture SYN_ARCH2 of ND2_611 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_610 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_610;

architecture SYN_ARCH2 of ND2_610 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_609 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_609;

architecture SYN_ARCH2 of ND2_609 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_608 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_608;

architecture SYN_ARCH2 of ND2_608 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_607 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_607;

architecture SYN_ARCH2 of ND2_607 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_606 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_606;

architecture SYN_ARCH2 of ND2_606 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_605 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_605;

architecture SYN_ARCH2 of ND2_605 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_604 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_604;

architecture SYN_ARCH2 of ND2_604 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_603 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_603;

architecture SYN_ARCH2 of ND2_603 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_602 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_602;

architecture SYN_ARCH2 of ND2_602 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_601 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_601;

architecture SYN_ARCH2 of ND2_601 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_600 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_600;

architecture SYN_ARCH2 of ND2_600 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_599 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_599;

architecture SYN_ARCH2 of ND2_599 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_598 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_598;

architecture SYN_ARCH2 of ND2_598 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_597 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_597;

architecture SYN_ARCH2 of ND2_597 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_596 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_596;

architecture SYN_ARCH2 of ND2_596 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_595 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_595;

architecture SYN_ARCH2 of ND2_595 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_594 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_594;

architecture SYN_ARCH2 of ND2_594 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_593 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_593;

architecture SYN_ARCH2 of ND2_593 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_592 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_592;

architecture SYN_ARCH2 of ND2_592 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_591 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_591;

architecture SYN_ARCH2 of ND2_591 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_590 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_590;

architecture SYN_ARCH2 of ND2_590 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_589 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_589;

architecture SYN_ARCH2 of ND2_589 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_588 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_588;

architecture SYN_ARCH2 of ND2_588 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_587 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_587;

architecture SYN_ARCH2 of ND2_587 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_586 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_586;

architecture SYN_ARCH2 of ND2_586 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_585 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_585;

architecture SYN_ARCH2 of ND2_585 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_584 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_584;

architecture SYN_ARCH2 of ND2_584 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_583 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_583;

architecture SYN_ARCH2 of ND2_583 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_582 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_582;

architecture SYN_ARCH2 of ND2_582 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_581 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_581;

architecture SYN_ARCH2 of ND2_581 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_580 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_580;

architecture SYN_ARCH2 of ND2_580 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_579 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_579;

architecture SYN_ARCH2 of ND2_579 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_578 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_578;

architecture SYN_ARCH2 of ND2_578 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_577 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_577;

architecture SYN_ARCH2 of ND2_577 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_576 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_576;

architecture SYN_ARCH2 of ND2_576 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_575 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_575;

architecture SYN_ARCH2 of ND2_575 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_574 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_574;

architecture SYN_ARCH2 of ND2_574 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_573 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_573;

architecture SYN_ARCH2 of ND2_573 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_572 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_572;

architecture SYN_ARCH2 of ND2_572 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_571 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_571;

architecture SYN_ARCH2 of ND2_571 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_570 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_570;

architecture SYN_ARCH2 of ND2_570 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_569 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_569;

architecture SYN_ARCH2 of ND2_569 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_568 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_568;

architecture SYN_ARCH2 of ND2_568 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_567 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_567;

architecture SYN_ARCH2 of ND2_567 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_566 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_566;

architecture SYN_ARCH2 of ND2_566 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_565 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_565;

architecture SYN_ARCH2 of ND2_565 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_564 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_564;

architecture SYN_ARCH2 of ND2_564 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_563 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_563;

architecture SYN_ARCH2 of ND2_563 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_562 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_562;

architecture SYN_ARCH2 of ND2_562 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_561 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_561;

architecture SYN_ARCH2 of ND2_561 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_560 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_560;

architecture SYN_ARCH2 of ND2_560 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_559 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_559;

architecture SYN_ARCH2 of ND2_559 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_558 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_558;

architecture SYN_ARCH2 of ND2_558 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_557 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_557;

architecture SYN_ARCH2 of ND2_557 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_556 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_556;

architecture SYN_ARCH2 of ND2_556 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_555 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_555;

architecture SYN_ARCH2 of ND2_555 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_554 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_554;

architecture SYN_ARCH2 of ND2_554 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_553 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_553;

architecture SYN_ARCH2 of ND2_553 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_552 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_552;

architecture SYN_ARCH2 of ND2_552 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_551 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_551;

architecture SYN_ARCH2 of ND2_551 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_550 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_550;

architecture SYN_ARCH2 of ND2_550 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_549 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_549;

architecture SYN_ARCH2 of ND2_549 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_548 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_548;

architecture SYN_ARCH2 of ND2_548 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_547 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_547;

architecture SYN_ARCH2 of ND2_547 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_546 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_546;

architecture SYN_ARCH2 of ND2_546 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_545 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_545;

architecture SYN_ARCH2 of ND2_545 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_544 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_544;

architecture SYN_ARCH2 of ND2_544 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_543 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_543;

architecture SYN_ARCH2 of ND2_543 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_542 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_542;

architecture SYN_ARCH2 of ND2_542 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_541 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_541;

architecture SYN_ARCH2 of ND2_541 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_540 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_540;

architecture SYN_ARCH2 of ND2_540 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_539 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_539;

architecture SYN_ARCH2 of ND2_539 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_538 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_538;

architecture SYN_ARCH2 of ND2_538 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_537 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_537;

architecture SYN_ARCH2 of ND2_537 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_536 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_536;

architecture SYN_ARCH2 of ND2_536 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_535 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_535;

architecture SYN_ARCH2 of ND2_535 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_534 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_534;

architecture SYN_ARCH2 of ND2_534 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_533 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_533;

architecture SYN_ARCH2 of ND2_533 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_532 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_532;

architecture SYN_ARCH2 of ND2_532 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_531 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_531;

architecture SYN_ARCH2 of ND2_531 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_530 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_530;

architecture SYN_ARCH2 of ND2_530 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_529 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_529;

architecture SYN_ARCH2 of ND2_529 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_528 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_528;

architecture SYN_ARCH2 of ND2_528 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_527 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_527;

architecture SYN_ARCH2 of ND2_527 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_526 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_526;

architecture SYN_ARCH2 of ND2_526 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_525 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_525;

architecture SYN_ARCH2 of ND2_525 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_524 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_524;

architecture SYN_ARCH2 of ND2_524 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_523 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_523;

architecture SYN_ARCH2 of ND2_523 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_522 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_522;

architecture SYN_ARCH2 of ND2_522 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_521 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_521;

architecture SYN_ARCH2 of ND2_521 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_520 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_520;

architecture SYN_ARCH2 of ND2_520 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_519 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_519;

architecture SYN_ARCH2 of ND2_519 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_518 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_518;

architecture SYN_ARCH2 of ND2_518 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_517 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_517;

architecture SYN_ARCH2 of ND2_517 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_516 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_516;

architecture SYN_ARCH2 of ND2_516 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_515 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_515;

architecture SYN_ARCH2 of ND2_515 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_514 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_514;

architecture SYN_ARCH2 of ND2_514 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_513 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_513;

architecture SYN_ARCH2 of ND2_513 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_512 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_512;

architecture SYN_ARCH2 of ND2_512 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_511 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_511;

architecture SYN_ARCH2 of ND2_511 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_510 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_510;

architecture SYN_ARCH2 of ND2_510 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_509 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_509;

architecture SYN_ARCH2 of ND2_509 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_508 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_508;

architecture SYN_ARCH2 of ND2_508 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_507 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_507;

architecture SYN_ARCH2 of ND2_507 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_506 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_506;

architecture SYN_ARCH2 of ND2_506 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_505 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_505;

architecture SYN_ARCH2 of ND2_505 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_504 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_504;

architecture SYN_ARCH2 of ND2_504 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_503 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_503;

architecture SYN_ARCH2 of ND2_503 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_502 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_502;

architecture SYN_ARCH2 of ND2_502 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_501 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_501;

architecture SYN_ARCH2 of ND2_501 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_500 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_500;

architecture SYN_ARCH2 of ND2_500 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_499 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_499;

architecture SYN_ARCH2 of ND2_499 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_498 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_498;

architecture SYN_ARCH2 of ND2_498 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_497 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_497;

architecture SYN_ARCH2 of ND2_497 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_496 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_496;

architecture SYN_ARCH2 of ND2_496 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_495 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_495;

architecture SYN_ARCH2 of ND2_495 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_494 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_494;

architecture SYN_ARCH2 of ND2_494 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_493 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_493;

architecture SYN_ARCH2 of ND2_493 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_492 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_492;

architecture SYN_ARCH2 of ND2_492 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_491 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_491;

architecture SYN_ARCH2 of ND2_491 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_490 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_490;

architecture SYN_ARCH2 of ND2_490 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_489 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_489;

architecture SYN_ARCH2 of ND2_489 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_488 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_488;

architecture SYN_ARCH2 of ND2_488 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_487 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_487;

architecture SYN_ARCH2 of ND2_487 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_486 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_486;

architecture SYN_ARCH2 of ND2_486 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_485 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_485;

architecture SYN_ARCH2 of ND2_485 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_484 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_484;

architecture SYN_ARCH2 of ND2_484 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_483 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_483;

architecture SYN_ARCH2 of ND2_483 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_482 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_482;

architecture SYN_ARCH2 of ND2_482 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_481 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_481;

architecture SYN_ARCH2 of ND2_481 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_480 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_480;

architecture SYN_ARCH2 of ND2_480 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_479 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_479;

architecture SYN_ARCH2 of ND2_479 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_478 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_478;

architecture SYN_ARCH2 of ND2_478 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_477 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_477;

architecture SYN_ARCH2 of ND2_477 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_476 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_476;

architecture SYN_ARCH2 of ND2_476 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_475 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_475;

architecture SYN_ARCH2 of ND2_475 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_474 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_474;

architecture SYN_ARCH2 of ND2_474 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_473 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_473;

architecture SYN_ARCH2 of ND2_473 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_472 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_472;

architecture SYN_ARCH2 of ND2_472 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_471 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_471;

architecture SYN_ARCH2 of ND2_471 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_470 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_470;

architecture SYN_ARCH2 of ND2_470 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_469 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_469;

architecture SYN_ARCH2 of ND2_469 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_468 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_468;

architecture SYN_ARCH2 of ND2_468 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_467 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_467;

architecture SYN_ARCH2 of ND2_467 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_466 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_466;

architecture SYN_ARCH2 of ND2_466 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_465 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_465;

architecture SYN_ARCH2 of ND2_465 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_464 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_464;

architecture SYN_ARCH2 of ND2_464 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_463 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_463;

architecture SYN_ARCH2 of ND2_463 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_462 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_462;

architecture SYN_ARCH2 of ND2_462 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_461 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_461;

architecture SYN_ARCH2 of ND2_461 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_460 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_460;

architecture SYN_ARCH2 of ND2_460 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_459 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_459;

architecture SYN_ARCH2 of ND2_459 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_458 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_458;

architecture SYN_ARCH2 of ND2_458 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_457 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_457;

architecture SYN_ARCH2 of ND2_457 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_456 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_456;

architecture SYN_ARCH2 of ND2_456 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_455 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_455;

architecture SYN_ARCH2 of ND2_455 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_454 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_454;

architecture SYN_ARCH2 of ND2_454 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_453 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_453;

architecture SYN_ARCH2 of ND2_453 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_452 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_452;

architecture SYN_ARCH2 of ND2_452 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_451 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_451;

architecture SYN_ARCH2 of ND2_451 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_450 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_450;

architecture SYN_ARCH2 of ND2_450 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_449 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_449;

architecture SYN_ARCH2 of ND2_449 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_448 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_448;

architecture SYN_ARCH2 of ND2_448 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_447 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_447;

architecture SYN_ARCH2 of ND2_447 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_446 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_446;

architecture SYN_ARCH2 of ND2_446 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_445 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_445;

architecture SYN_ARCH2 of ND2_445 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_444 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_444;

architecture SYN_ARCH2 of ND2_444 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_443 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_443;

architecture SYN_ARCH2 of ND2_443 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_442 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_442;

architecture SYN_ARCH2 of ND2_442 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_441 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_441;

architecture SYN_ARCH2 of ND2_441 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_440 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_440;

architecture SYN_ARCH2 of ND2_440 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_439 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_439;

architecture SYN_ARCH2 of ND2_439 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_438 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_438;

architecture SYN_ARCH2 of ND2_438 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_437 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_437;

architecture SYN_ARCH2 of ND2_437 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_436 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_436;

architecture SYN_ARCH2 of ND2_436 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_435 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_435;

architecture SYN_ARCH2 of ND2_435 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_434 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_434;

architecture SYN_ARCH2 of ND2_434 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_433 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_433;

architecture SYN_ARCH2 of ND2_433 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_432 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_432;

architecture SYN_ARCH2 of ND2_432 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_431 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_431;

architecture SYN_ARCH2 of ND2_431 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_430 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_430;

architecture SYN_ARCH2 of ND2_430 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_429 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_429;

architecture SYN_ARCH2 of ND2_429 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_428 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_428;

architecture SYN_ARCH2 of ND2_428 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_427 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_427;

architecture SYN_ARCH2 of ND2_427 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_426 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_426;

architecture SYN_ARCH2 of ND2_426 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_425 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_425;

architecture SYN_ARCH2 of ND2_425 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_424 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_424;

architecture SYN_ARCH2 of ND2_424 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_423 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_423;

architecture SYN_ARCH2 of ND2_423 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_422 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_422;

architecture SYN_ARCH2 of ND2_422 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_421 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_421;

architecture SYN_ARCH2 of ND2_421 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_420 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_420;

architecture SYN_ARCH2 of ND2_420 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_419 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_419;

architecture SYN_ARCH2 of ND2_419 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_418 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_418;

architecture SYN_ARCH2 of ND2_418 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_417 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_417;

architecture SYN_ARCH2 of ND2_417 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_416 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_416;

architecture SYN_ARCH2 of ND2_416 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_415 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_415;

architecture SYN_ARCH2 of ND2_415 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_414 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_414;

architecture SYN_ARCH2 of ND2_414 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_413 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_413;

architecture SYN_ARCH2 of ND2_413 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_412 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_412;

architecture SYN_ARCH2 of ND2_412 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_411 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_411;

architecture SYN_ARCH2 of ND2_411 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_410 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_410;

architecture SYN_ARCH2 of ND2_410 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_409 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_409;

architecture SYN_ARCH2 of ND2_409 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_408 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_408;

architecture SYN_ARCH2 of ND2_408 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_407 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_407;

architecture SYN_ARCH2 of ND2_407 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_406 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_406;

architecture SYN_ARCH2 of ND2_406 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_405 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_405;

architecture SYN_ARCH2 of ND2_405 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_404 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_404;

architecture SYN_ARCH2 of ND2_404 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_403 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_403;

architecture SYN_ARCH2 of ND2_403 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_402 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_402;

architecture SYN_ARCH2 of ND2_402 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_401 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_401;

architecture SYN_ARCH2 of ND2_401 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_400 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_400;

architecture SYN_ARCH2 of ND2_400 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_399 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_399;

architecture SYN_ARCH2 of ND2_399 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_398 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_398;

architecture SYN_ARCH2 of ND2_398 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_397 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_397;

architecture SYN_ARCH2 of ND2_397 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_396 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_396;

architecture SYN_ARCH2 of ND2_396 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_395 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_395;

architecture SYN_ARCH2 of ND2_395 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_394 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_394;

architecture SYN_ARCH2 of ND2_394 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_393 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_393;

architecture SYN_ARCH2 of ND2_393 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_392 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_392;

architecture SYN_ARCH2 of ND2_392 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_391 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_391;

architecture SYN_ARCH2 of ND2_391 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_390 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_390;

architecture SYN_ARCH2 of ND2_390 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_389 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_389;

architecture SYN_ARCH2 of ND2_389 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_388 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_388;

architecture SYN_ARCH2 of ND2_388 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_387 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_387;

architecture SYN_ARCH2 of ND2_387 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_386 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_386;

architecture SYN_ARCH2 of ND2_386 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_385 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_385;

architecture SYN_ARCH2 of ND2_385 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_384 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_384;

architecture SYN_ARCH2 of ND2_384 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_383 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_383;

architecture SYN_ARCH2 of ND2_383 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_382 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_382;

architecture SYN_ARCH2 of ND2_382 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_381 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_381;

architecture SYN_ARCH2 of ND2_381 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_380 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_380;

architecture SYN_ARCH2 of ND2_380 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_379 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_379;

architecture SYN_ARCH2 of ND2_379 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_378 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_378;

architecture SYN_ARCH2 of ND2_378 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_377 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_377;

architecture SYN_ARCH2 of ND2_377 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_376 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_376;

architecture SYN_ARCH2 of ND2_376 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_375 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_375;

architecture SYN_ARCH2 of ND2_375 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_374 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_374;

architecture SYN_ARCH2 of ND2_374 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_373 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_373;

architecture SYN_ARCH2 of ND2_373 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_372 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_372;

architecture SYN_ARCH2 of ND2_372 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_371 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_371;

architecture SYN_ARCH2 of ND2_371 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_370 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_370;

architecture SYN_ARCH2 of ND2_370 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_369 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_369;

architecture SYN_ARCH2 of ND2_369 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_368 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_368;

architecture SYN_ARCH2 of ND2_368 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_367 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_367;

architecture SYN_ARCH2 of ND2_367 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_366 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_366;

architecture SYN_ARCH2 of ND2_366 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_365 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_365;

architecture SYN_ARCH2 of ND2_365 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_364 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_364;

architecture SYN_ARCH2 of ND2_364 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_363 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_363;

architecture SYN_ARCH2 of ND2_363 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_362 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_362;

architecture SYN_ARCH2 of ND2_362 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_361 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_361;

architecture SYN_ARCH2 of ND2_361 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_360 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_360;

architecture SYN_ARCH2 of ND2_360 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_359 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_359;

architecture SYN_ARCH2 of ND2_359 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_358 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_358;

architecture SYN_ARCH2 of ND2_358 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_357 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_357;

architecture SYN_ARCH2 of ND2_357 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_356 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_356;

architecture SYN_ARCH2 of ND2_356 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_355 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_355;

architecture SYN_ARCH2 of ND2_355 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_354 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_354;

architecture SYN_ARCH2 of ND2_354 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_353 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_353;

architecture SYN_ARCH2 of ND2_353 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_352 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_352;

architecture SYN_ARCH2 of ND2_352 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_351 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_351;

architecture SYN_ARCH2 of ND2_351 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_350 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_350;

architecture SYN_ARCH2 of ND2_350 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_349 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_349;

architecture SYN_ARCH2 of ND2_349 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_348 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_348;

architecture SYN_ARCH2 of ND2_348 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_347 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_347;

architecture SYN_ARCH2 of ND2_347 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_346 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_346;

architecture SYN_ARCH2 of ND2_346 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_345 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_345;

architecture SYN_ARCH2 of ND2_345 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_344 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_344;

architecture SYN_ARCH2 of ND2_344 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_343 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_343;

architecture SYN_ARCH2 of ND2_343 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_342 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_342;

architecture SYN_ARCH2 of ND2_342 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_341 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_341;

architecture SYN_ARCH2 of ND2_341 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_340 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_340;

architecture SYN_ARCH2 of ND2_340 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_339 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_339;

architecture SYN_ARCH2 of ND2_339 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_338 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_338;

architecture SYN_ARCH2 of ND2_338 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_337 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_337;

architecture SYN_ARCH2 of ND2_337 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_336 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_336;

architecture SYN_ARCH2 of ND2_336 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_335 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_335;

architecture SYN_ARCH2 of ND2_335 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_334 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_334;

architecture SYN_ARCH2 of ND2_334 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_333 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_333;

architecture SYN_ARCH2 of ND2_333 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_332 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_332;

architecture SYN_ARCH2 of ND2_332 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_331 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_331;

architecture SYN_ARCH2 of ND2_331 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_330 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_330;

architecture SYN_ARCH2 of ND2_330 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_329 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_329;

architecture SYN_ARCH2 of ND2_329 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_328 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_328;

architecture SYN_ARCH2 of ND2_328 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_327 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_327;

architecture SYN_ARCH2 of ND2_327 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_326 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_326;

architecture SYN_ARCH2 of ND2_326 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_325 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_325;

architecture SYN_ARCH2 of ND2_325 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_324 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_324;

architecture SYN_ARCH2 of ND2_324 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_323 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_323;

architecture SYN_ARCH2 of ND2_323 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_322 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_322;

architecture SYN_ARCH2 of ND2_322 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_321 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_321;

architecture SYN_ARCH2 of ND2_321 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_320 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_320;

architecture SYN_ARCH2 of ND2_320 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_319 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_319;

architecture SYN_ARCH2 of ND2_319 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_318 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_318;

architecture SYN_ARCH2 of ND2_318 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_317 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_317;

architecture SYN_ARCH2 of ND2_317 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_316 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_316;

architecture SYN_ARCH2 of ND2_316 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_315 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_315;

architecture SYN_ARCH2 of ND2_315 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_314 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_314;

architecture SYN_ARCH2 of ND2_314 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_313 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_313;

architecture SYN_ARCH2 of ND2_313 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_312 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_312;

architecture SYN_ARCH2 of ND2_312 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_311 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_311;

architecture SYN_ARCH2 of ND2_311 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_310 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_310;

architecture SYN_ARCH2 of ND2_310 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_309 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_309;

architecture SYN_ARCH2 of ND2_309 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_308 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_308;

architecture SYN_ARCH2 of ND2_308 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_307 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_307;

architecture SYN_ARCH2 of ND2_307 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_306 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_306;

architecture SYN_ARCH2 of ND2_306 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_305 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_305;

architecture SYN_ARCH2 of ND2_305 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_304 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_304;

architecture SYN_ARCH2 of ND2_304 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_303 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_303;

architecture SYN_ARCH2 of ND2_303 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_302 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_302;

architecture SYN_ARCH2 of ND2_302 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_301 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_301;

architecture SYN_ARCH2 of ND2_301 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_300 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_300;

architecture SYN_ARCH2 of ND2_300 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_299 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_299;

architecture SYN_ARCH2 of ND2_299 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_298 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_298;

architecture SYN_ARCH2 of ND2_298 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_297 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_297;

architecture SYN_ARCH2 of ND2_297 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_296 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_296;

architecture SYN_ARCH2 of ND2_296 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_295 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_295;

architecture SYN_ARCH2 of ND2_295 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_294 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_294;

architecture SYN_ARCH2 of ND2_294 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_293 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_293;

architecture SYN_ARCH2 of ND2_293 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_292 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_292;

architecture SYN_ARCH2 of ND2_292 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_291 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_291;

architecture SYN_ARCH2 of ND2_291 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_290 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_290;

architecture SYN_ARCH2 of ND2_290 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_289 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_289;

architecture SYN_ARCH2 of ND2_289 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_288 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_288;

architecture SYN_ARCH2 of ND2_288 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_287 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_287;

architecture SYN_ARCH2 of ND2_287 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_286 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_286;

architecture SYN_ARCH2 of ND2_286 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_285 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_285;

architecture SYN_ARCH2 of ND2_285 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_284 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_284;

architecture SYN_ARCH2 of ND2_284 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_283 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_283;

architecture SYN_ARCH2 of ND2_283 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_282 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_282;

architecture SYN_ARCH2 of ND2_282 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_281 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_281;

architecture SYN_ARCH2 of ND2_281 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_280 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_280;

architecture SYN_ARCH2 of ND2_280 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_279 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_279;

architecture SYN_ARCH2 of ND2_279 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_278 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_278;

architecture SYN_ARCH2 of ND2_278 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_277 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_277;

architecture SYN_ARCH2 of ND2_277 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_276 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_276;

architecture SYN_ARCH2 of ND2_276 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_275 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_275;

architecture SYN_ARCH2 of ND2_275 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_274 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_274;

architecture SYN_ARCH2 of ND2_274 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_273 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_273;

architecture SYN_ARCH2 of ND2_273 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_272 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_272;

architecture SYN_ARCH2 of ND2_272 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_271 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_271;

architecture SYN_ARCH2 of ND2_271 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_270 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_270;

architecture SYN_ARCH2 of ND2_270 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_269 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_269;

architecture SYN_ARCH2 of ND2_269 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_268 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_268;

architecture SYN_ARCH2 of ND2_268 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_267 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_267;

architecture SYN_ARCH2 of ND2_267 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_266 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_266;

architecture SYN_ARCH2 of ND2_266 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_265 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_265;

architecture SYN_ARCH2 of ND2_265 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_264 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_264;

architecture SYN_ARCH2 of ND2_264 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_263 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_263;

architecture SYN_ARCH2 of ND2_263 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_262 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_262;

architecture SYN_ARCH2 of ND2_262 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_261 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_261;

architecture SYN_ARCH2 of ND2_261 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_260 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_260;

architecture SYN_ARCH2 of ND2_260 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_259 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_259;

architecture SYN_ARCH2 of ND2_259 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_258 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_258;

architecture SYN_ARCH2 of ND2_258 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_257 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_257;

architecture SYN_ARCH2 of ND2_257 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_256 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_256;

architecture SYN_ARCH2 of ND2_256 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_255 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_255;

architecture SYN_ARCH2 of ND2_255 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_254 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_254;

architecture SYN_ARCH2 of ND2_254 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_253 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_253;

architecture SYN_ARCH2 of ND2_253 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_252 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_252;

architecture SYN_ARCH2 of ND2_252 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_251 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_251;

architecture SYN_ARCH2 of ND2_251 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_250 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_250;

architecture SYN_ARCH2 of ND2_250 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_249 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_249;

architecture SYN_ARCH2 of ND2_249 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_248 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_248;

architecture SYN_ARCH2 of ND2_248 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_247 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_247;

architecture SYN_ARCH2 of ND2_247 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_246 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_246;

architecture SYN_ARCH2 of ND2_246 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_245 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_245;

architecture SYN_ARCH2 of ND2_245 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_244 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_244;

architecture SYN_ARCH2 of ND2_244 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_243 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_243;

architecture SYN_ARCH2 of ND2_243 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_242 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_242;

architecture SYN_ARCH2 of ND2_242 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_241 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_241;

architecture SYN_ARCH2 of ND2_241 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_240 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_240;

architecture SYN_ARCH2 of ND2_240 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_239 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_239;

architecture SYN_ARCH2 of ND2_239 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_238 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_238;

architecture SYN_ARCH2 of ND2_238 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_237 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_237;

architecture SYN_ARCH2 of ND2_237 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_236 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_236;

architecture SYN_ARCH2 of ND2_236 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_235 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_235;

architecture SYN_ARCH2 of ND2_235 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_234 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_234;

architecture SYN_ARCH2 of ND2_234 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_233 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_233;

architecture SYN_ARCH2 of ND2_233 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_232 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_232;

architecture SYN_ARCH2 of ND2_232 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_231 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_231;

architecture SYN_ARCH2 of ND2_231 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_230 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_230;

architecture SYN_ARCH2 of ND2_230 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_229 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_229;

architecture SYN_ARCH2 of ND2_229 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_228 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_228;

architecture SYN_ARCH2 of ND2_228 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_227 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_227;

architecture SYN_ARCH2 of ND2_227 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_226 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_226;

architecture SYN_ARCH2 of ND2_226 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_225 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_225;

architecture SYN_ARCH2 of ND2_225 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_224 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_224;

architecture SYN_ARCH2 of ND2_224 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_223 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_223;

architecture SYN_ARCH2 of ND2_223 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_222 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_222;

architecture SYN_ARCH2 of ND2_222 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_221 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_221;

architecture SYN_ARCH2 of ND2_221 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_220 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_220;

architecture SYN_ARCH2 of ND2_220 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_219 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_219;

architecture SYN_ARCH2 of ND2_219 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_218 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_218;

architecture SYN_ARCH2 of ND2_218 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_217 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_217;

architecture SYN_ARCH2 of ND2_217 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_216 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_216;

architecture SYN_ARCH2 of ND2_216 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_215 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_215;

architecture SYN_ARCH2 of ND2_215 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_214 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_214;

architecture SYN_ARCH2 of ND2_214 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_213 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_213;

architecture SYN_ARCH2 of ND2_213 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_212 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_212;

architecture SYN_ARCH2 of ND2_212 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_211 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_211;

architecture SYN_ARCH2 of ND2_211 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_210 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_210;

architecture SYN_ARCH2 of ND2_210 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_209 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_209;

architecture SYN_ARCH2 of ND2_209 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_208 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_208;

architecture SYN_ARCH2 of ND2_208 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_207 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_207;

architecture SYN_ARCH2 of ND2_207 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_206 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_206;

architecture SYN_ARCH2 of ND2_206 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_205 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_205;

architecture SYN_ARCH2 of ND2_205 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_204 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_204;

architecture SYN_ARCH2 of ND2_204 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_203 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_203;

architecture SYN_ARCH2 of ND2_203 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_202 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_202;

architecture SYN_ARCH2 of ND2_202 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_201 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_201;

architecture SYN_ARCH2 of ND2_201 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_200 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_200;

architecture SYN_ARCH2 of ND2_200 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_199 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_199;

architecture SYN_ARCH2 of ND2_199 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_198 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_198;

architecture SYN_ARCH2 of ND2_198 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_197 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_197;

architecture SYN_ARCH2 of ND2_197 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_196 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_196;

architecture SYN_ARCH2 of ND2_196 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_195 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_195;

architecture SYN_ARCH2 of ND2_195 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_194 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_194;

architecture SYN_ARCH2 of ND2_194 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_193 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_193;

architecture SYN_ARCH2 of ND2_193 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_192 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_192;

architecture SYN_ARCH2 of ND2_192 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_191 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_191;

architecture SYN_ARCH2 of ND2_191 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_190 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_190;

architecture SYN_ARCH2 of ND2_190 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_189 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_189;

architecture SYN_ARCH2 of ND2_189 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_188 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_188;

architecture SYN_ARCH2 of ND2_188 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_187 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_187;

architecture SYN_ARCH2 of ND2_187 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_186 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_186;

architecture SYN_ARCH2 of ND2_186 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_185 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_185;

architecture SYN_ARCH2 of ND2_185 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_184 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_184;

architecture SYN_ARCH2 of ND2_184 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_183 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_183;

architecture SYN_ARCH2 of ND2_183 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_182 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_182;

architecture SYN_ARCH2 of ND2_182 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_181 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_181;

architecture SYN_ARCH2 of ND2_181 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_180 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_180;

architecture SYN_ARCH2 of ND2_180 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_179 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_179;

architecture SYN_ARCH2 of ND2_179 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_178 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_178;

architecture SYN_ARCH2 of ND2_178 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_177 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_177;

architecture SYN_ARCH2 of ND2_177 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_176 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_176;

architecture SYN_ARCH2 of ND2_176 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_175 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_175;

architecture SYN_ARCH2 of ND2_175 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_174 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_174;

architecture SYN_ARCH2 of ND2_174 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_173 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_173;

architecture SYN_ARCH2 of ND2_173 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_172 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_172;

architecture SYN_ARCH2 of ND2_172 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_171 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_171;

architecture SYN_ARCH2 of ND2_171 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_170 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_170;

architecture SYN_ARCH2 of ND2_170 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_169 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_169;

architecture SYN_ARCH2 of ND2_169 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_168 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_168;

architecture SYN_ARCH2 of ND2_168 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_167 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_167;

architecture SYN_ARCH2 of ND2_167 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_166 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_166;

architecture SYN_ARCH2 of ND2_166 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_165 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_165;

architecture SYN_ARCH2 of ND2_165 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_164 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_164;

architecture SYN_ARCH2 of ND2_164 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_163 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_163;

architecture SYN_ARCH2 of ND2_163 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_162 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_162;

architecture SYN_ARCH2 of ND2_162 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_161 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_161;

architecture SYN_ARCH2 of ND2_161 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_160 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_160;

architecture SYN_ARCH2 of ND2_160 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_159 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_159;

architecture SYN_ARCH2 of ND2_159 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_158 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_158;

architecture SYN_ARCH2 of ND2_158 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_157 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_157;

architecture SYN_ARCH2 of ND2_157 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_156 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_156;

architecture SYN_ARCH2 of ND2_156 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_155 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_155;

architecture SYN_ARCH2 of ND2_155 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_154 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_154;

architecture SYN_ARCH2 of ND2_154 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_153 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_153;

architecture SYN_ARCH2 of ND2_153 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_152 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_152;

architecture SYN_ARCH2 of ND2_152 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_151 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_151;

architecture SYN_ARCH2 of ND2_151 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_150 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_150;

architecture SYN_ARCH2 of ND2_150 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_149 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_149;

architecture SYN_ARCH2 of ND2_149 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_148 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_148;

architecture SYN_ARCH2 of ND2_148 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_147 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_147;

architecture SYN_ARCH2 of ND2_147 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_146 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_146;

architecture SYN_ARCH2 of ND2_146 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_145 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_145;

architecture SYN_ARCH2 of ND2_145 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_144 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_144;

architecture SYN_ARCH2 of ND2_144 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_143 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_143;

architecture SYN_ARCH2 of ND2_143 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_142 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_142;

architecture SYN_ARCH2 of ND2_142 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_141 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_141;

architecture SYN_ARCH2 of ND2_141 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_140 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_140;

architecture SYN_ARCH2 of ND2_140 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_139 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_139;

architecture SYN_ARCH2 of ND2_139 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_138 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_138;

architecture SYN_ARCH2 of ND2_138 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_137 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_137;

architecture SYN_ARCH2 of ND2_137 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_136 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_136;

architecture SYN_ARCH2 of ND2_136 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_135 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_135;

architecture SYN_ARCH2 of ND2_135 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_134 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_134;

architecture SYN_ARCH2 of ND2_134 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_133 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_133;

architecture SYN_ARCH2 of ND2_133 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_132 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_132;

architecture SYN_ARCH2 of ND2_132 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_131 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_131;

architecture SYN_ARCH2 of ND2_131 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_130 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_130;

architecture SYN_ARCH2 of ND2_130 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_129 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_129;

architecture SYN_ARCH2 of ND2_129 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_128 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_128;

architecture SYN_ARCH2 of ND2_128 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_127 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_127;

architecture SYN_ARCH2 of ND2_127 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_126 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_126;

architecture SYN_ARCH2 of ND2_126 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_125 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_125;

architecture SYN_ARCH2 of ND2_125 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_124 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_124;

architecture SYN_ARCH2 of ND2_124 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_123 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_123;

architecture SYN_ARCH2 of ND2_123 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_122 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_122;

architecture SYN_ARCH2 of ND2_122 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_121 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_121;

architecture SYN_ARCH2 of ND2_121 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_120 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_120;

architecture SYN_ARCH2 of ND2_120 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_119 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_119;

architecture SYN_ARCH2 of ND2_119 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_118 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_118;

architecture SYN_ARCH2 of ND2_118 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_117 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_117;

architecture SYN_ARCH2 of ND2_117 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_116 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_116;

architecture SYN_ARCH2 of ND2_116 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_115 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_115;

architecture SYN_ARCH2 of ND2_115 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_114 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_114;

architecture SYN_ARCH2 of ND2_114 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_113 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_113;

architecture SYN_ARCH2 of ND2_113 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_112 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_112;

architecture SYN_ARCH2 of ND2_112 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_111 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_111;

architecture SYN_ARCH2 of ND2_111 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_110 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_110;

architecture SYN_ARCH2 of ND2_110 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_109 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_109;

architecture SYN_ARCH2 of ND2_109 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_108 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_108;

architecture SYN_ARCH2 of ND2_108 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_107 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_107;

architecture SYN_ARCH2 of ND2_107 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_106 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_106;

architecture SYN_ARCH2 of ND2_106 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_105 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_105;

architecture SYN_ARCH2 of ND2_105 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_104 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_104;

architecture SYN_ARCH2 of ND2_104 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_103 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_103;

architecture SYN_ARCH2 of ND2_103 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_102 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_102;

architecture SYN_ARCH2 of ND2_102 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_101 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_101;

architecture SYN_ARCH2 of ND2_101 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_100 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_100;

architecture SYN_ARCH2 of ND2_100 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_99 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_99;

architecture SYN_ARCH2 of ND2_99 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_98 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_98;

architecture SYN_ARCH2 of ND2_98 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_97 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_97;

architecture SYN_ARCH2 of ND2_97 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_96 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_96;

architecture SYN_ARCH2 of ND2_96 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_95 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_95;

architecture SYN_ARCH2 of ND2_95 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_94 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_94;

architecture SYN_ARCH2 of ND2_94 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_93 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_93;

architecture SYN_ARCH2 of ND2_93 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_92 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_92;

architecture SYN_ARCH2 of ND2_92 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_91 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_91;

architecture SYN_ARCH2 of ND2_91 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_90 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_90;

architecture SYN_ARCH2 of ND2_90 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_89 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_89;

architecture SYN_ARCH2 of ND2_89 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_88 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_88;

architecture SYN_ARCH2 of ND2_88 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_87 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_87;

architecture SYN_ARCH2 of ND2_87 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_86 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_86;

architecture SYN_ARCH2 of ND2_86 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_85 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_85;

architecture SYN_ARCH2 of ND2_85 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_84 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_84;

architecture SYN_ARCH2 of ND2_84 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_83 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_83;

architecture SYN_ARCH2 of ND2_83 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_82 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_82;

architecture SYN_ARCH2 of ND2_82 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_81 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_81;

architecture SYN_ARCH2 of ND2_81 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_80 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_80;

architecture SYN_ARCH2 of ND2_80 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_79 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_79;

architecture SYN_ARCH2 of ND2_79 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_78 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_78;

architecture SYN_ARCH2 of ND2_78 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_77 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_77;

architecture SYN_ARCH2 of ND2_77 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_76 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_76;

architecture SYN_ARCH2 of ND2_76 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_75 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_75;

architecture SYN_ARCH2 of ND2_75 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_74 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_74;

architecture SYN_ARCH2 of ND2_74 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_73 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_73;

architecture SYN_ARCH2 of ND2_73 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_72 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_72;

architecture SYN_ARCH2 of ND2_72 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_71 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_71;

architecture SYN_ARCH2 of ND2_71 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_70 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_70;

architecture SYN_ARCH2 of ND2_70 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_69 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_69;

architecture SYN_ARCH2 of ND2_69 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_68 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_68;

architecture SYN_ARCH2 of ND2_68 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_67 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_67;

architecture SYN_ARCH2 of ND2_67 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_66 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_66;

architecture SYN_ARCH2 of ND2_66 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_65 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_65;

architecture SYN_ARCH2 of ND2_65 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_64 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_64;

architecture SYN_ARCH2 of ND2_64 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_63 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_63;

architecture SYN_ARCH2 of ND2_63 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_62 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_62;

architecture SYN_ARCH2 of ND2_62 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_61 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_61;

architecture SYN_ARCH2 of ND2_61 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_60 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_60;

architecture SYN_ARCH2 of ND2_60 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_59 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_59;

architecture SYN_ARCH2 of ND2_59 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_58 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_58;

architecture SYN_ARCH2 of ND2_58 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_57 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_57;

architecture SYN_ARCH2 of ND2_57 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_56 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_56;

architecture SYN_ARCH2 of ND2_56 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_55 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_55;

architecture SYN_ARCH2 of ND2_55 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_54 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_54;

architecture SYN_ARCH2 of ND2_54 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_53 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_53;

architecture SYN_ARCH2 of ND2_53 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_52 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_52;

architecture SYN_ARCH2 of ND2_52 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_51 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_51;

architecture SYN_ARCH2 of ND2_51 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_50 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_50;

architecture SYN_ARCH2 of ND2_50 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_49 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_49;

architecture SYN_ARCH2 of ND2_49 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_48 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_48;

architecture SYN_ARCH2 of ND2_48 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_47 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_47;

architecture SYN_ARCH2 of ND2_47 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_46 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_46;

architecture SYN_ARCH2 of ND2_46 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_45 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_45;

architecture SYN_ARCH2 of ND2_45 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_44 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_44;

architecture SYN_ARCH2 of ND2_44 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_43 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_43;

architecture SYN_ARCH2 of ND2_43 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_42 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_42;

architecture SYN_ARCH2 of ND2_42 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_41 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_41;

architecture SYN_ARCH2 of ND2_41 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_40 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_40;

architecture SYN_ARCH2 of ND2_40 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_39 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_39;

architecture SYN_ARCH2 of ND2_39 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_38 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_38;

architecture SYN_ARCH2 of ND2_38 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_37 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_37;

architecture SYN_ARCH2 of ND2_37 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_36 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_36;

architecture SYN_ARCH2 of ND2_36 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_35 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_35;

architecture SYN_ARCH2 of ND2_35 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_34 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_34;

architecture SYN_ARCH2 of ND2_34 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_33 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_33;

architecture SYN_ARCH2 of ND2_33 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_32 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_32;

architecture SYN_ARCH2 of ND2_32 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_31 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_31;

architecture SYN_ARCH2 of ND2_31 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_30 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_30;

architecture SYN_ARCH2 of ND2_30 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_29 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_29;

architecture SYN_ARCH2 of ND2_29 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_28 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_28;

architecture SYN_ARCH2 of ND2_28 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_27 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_27;

architecture SYN_ARCH2 of ND2_27 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_26 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_26;

architecture SYN_ARCH2 of ND2_26 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_25 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_25;

architecture SYN_ARCH2 of ND2_25 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_24 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_24;

architecture SYN_ARCH2 of ND2_24 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_23 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_23;

architecture SYN_ARCH2 of ND2_23 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_22 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_22;

architecture SYN_ARCH2 of ND2_22 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_21 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_21;

architecture SYN_ARCH2 of ND2_21 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_20 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_20;

architecture SYN_ARCH2 of ND2_20 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_19 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_19;

architecture SYN_ARCH2 of ND2_19 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_18 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_18;

architecture SYN_ARCH2 of ND2_18 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_17 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_17;

architecture SYN_ARCH2 of ND2_17 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_16 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_16;

architecture SYN_ARCH2 of ND2_16 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_15 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_15;

architecture SYN_ARCH2 of ND2_15 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_14 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_14;

architecture SYN_ARCH2 of ND2_14 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_13 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_13;

architecture SYN_ARCH2 of ND2_13 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_12 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_12;

architecture SYN_ARCH2 of ND2_12 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_11 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_11;

architecture SYN_ARCH2 of ND2_11 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_10 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_10;

architecture SYN_ARCH2 of ND2_10 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_9 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_9;

architecture SYN_ARCH2 of ND2_9 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_8 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_8;

architecture SYN_ARCH2 of ND2_8 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_7 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_7;

architecture SYN_ARCH2 of ND2_7 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_6 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_6;

architecture SYN_ARCH2 of ND2_6 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_5 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_5;

architecture SYN_ARCH2 of ND2_5 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_4 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_4;

architecture SYN_ARCH2 of ND2_4 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_3 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_3;

architecture SYN_ARCH2 of ND2_3 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_2 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_2;

architecture SYN_ARCH2 of ND2_2 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_1 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_1;

architecture SYN_ARCH2 of ND2_1 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_255 is

   port( A : in std_logic;  Y : out std_logic);

end IV_255;

architecture SYN_BEHAVIORAL of IV_255 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_254 is

   port( A : in std_logic;  Y : out std_logic);

end IV_254;

architecture SYN_BEHAVIORAL of IV_254 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_253 is

   port( A : in std_logic;  Y : out std_logic);

end IV_253;

architecture SYN_BEHAVIORAL of IV_253 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_252 is

   port( A : in std_logic;  Y : out std_logic);

end IV_252;

architecture SYN_BEHAVIORAL of IV_252 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_251 is

   port( A : in std_logic;  Y : out std_logic);

end IV_251;

architecture SYN_BEHAVIORAL of IV_251 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_250 is

   port( A : in std_logic;  Y : out std_logic);

end IV_250;

architecture SYN_BEHAVIORAL of IV_250 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_249 is

   port( A : in std_logic;  Y : out std_logic);

end IV_249;

architecture SYN_BEHAVIORAL of IV_249 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_248 is

   port( A : in std_logic;  Y : out std_logic);

end IV_248;

architecture SYN_BEHAVIORAL of IV_248 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_247 is

   port( A : in std_logic;  Y : out std_logic);

end IV_247;

architecture SYN_BEHAVIORAL of IV_247 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_246 is

   port( A : in std_logic;  Y : out std_logic);

end IV_246;

architecture SYN_BEHAVIORAL of IV_246 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_245 is

   port( A : in std_logic;  Y : out std_logic);

end IV_245;

architecture SYN_BEHAVIORAL of IV_245 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_244 is

   port( A : in std_logic;  Y : out std_logic);

end IV_244;

architecture SYN_BEHAVIORAL of IV_244 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_243 is

   port( A : in std_logic;  Y : out std_logic);

end IV_243;

architecture SYN_BEHAVIORAL of IV_243 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_242 is

   port( A : in std_logic;  Y : out std_logic);

end IV_242;

architecture SYN_BEHAVIORAL of IV_242 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_241 is

   port( A : in std_logic;  Y : out std_logic);

end IV_241;

architecture SYN_BEHAVIORAL of IV_241 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_240 is

   port( A : in std_logic;  Y : out std_logic);

end IV_240;

architecture SYN_BEHAVIORAL of IV_240 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_239 is

   port( A : in std_logic;  Y : out std_logic);

end IV_239;

architecture SYN_BEHAVIORAL of IV_239 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_238 is

   port( A : in std_logic;  Y : out std_logic);

end IV_238;

architecture SYN_BEHAVIORAL of IV_238 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_237 is

   port( A : in std_logic;  Y : out std_logic);

end IV_237;

architecture SYN_BEHAVIORAL of IV_237 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_236 is

   port( A : in std_logic;  Y : out std_logic);

end IV_236;

architecture SYN_BEHAVIORAL of IV_236 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_235 is

   port( A : in std_logic;  Y : out std_logic);

end IV_235;

architecture SYN_BEHAVIORAL of IV_235 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_234 is

   port( A : in std_logic;  Y : out std_logic);

end IV_234;

architecture SYN_BEHAVIORAL of IV_234 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_233 is

   port( A : in std_logic;  Y : out std_logic);

end IV_233;

architecture SYN_BEHAVIORAL of IV_233 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_232 is

   port( A : in std_logic;  Y : out std_logic);

end IV_232;

architecture SYN_BEHAVIORAL of IV_232 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_231 is

   port( A : in std_logic;  Y : out std_logic);

end IV_231;

architecture SYN_BEHAVIORAL of IV_231 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_230 is

   port( A : in std_logic;  Y : out std_logic);

end IV_230;

architecture SYN_BEHAVIORAL of IV_230 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_229 is

   port( A : in std_logic;  Y : out std_logic);

end IV_229;

architecture SYN_BEHAVIORAL of IV_229 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_228 is

   port( A : in std_logic;  Y : out std_logic);

end IV_228;

architecture SYN_BEHAVIORAL of IV_228 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_227 is

   port( A : in std_logic;  Y : out std_logic);

end IV_227;

architecture SYN_BEHAVIORAL of IV_227 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_226 is

   port( A : in std_logic;  Y : out std_logic);

end IV_226;

architecture SYN_BEHAVIORAL of IV_226 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_225 is

   port( A : in std_logic;  Y : out std_logic);

end IV_225;

architecture SYN_BEHAVIORAL of IV_225 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_224 is

   port( A : in std_logic;  Y : out std_logic);

end IV_224;

architecture SYN_BEHAVIORAL of IV_224 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_223 is

   port( A : in std_logic;  Y : out std_logic);

end IV_223;

architecture SYN_BEHAVIORAL of IV_223 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_222 is

   port( A : in std_logic;  Y : out std_logic);

end IV_222;

architecture SYN_BEHAVIORAL of IV_222 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_221 is

   port( A : in std_logic;  Y : out std_logic);

end IV_221;

architecture SYN_BEHAVIORAL of IV_221 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_220 is

   port( A : in std_logic;  Y : out std_logic);

end IV_220;

architecture SYN_BEHAVIORAL of IV_220 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_219 is

   port( A : in std_logic;  Y : out std_logic);

end IV_219;

architecture SYN_BEHAVIORAL of IV_219 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_218 is

   port( A : in std_logic;  Y : out std_logic);

end IV_218;

architecture SYN_BEHAVIORAL of IV_218 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_217 is

   port( A : in std_logic;  Y : out std_logic);

end IV_217;

architecture SYN_BEHAVIORAL of IV_217 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_216 is

   port( A : in std_logic;  Y : out std_logic);

end IV_216;

architecture SYN_BEHAVIORAL of IV_216 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_215 is

   port( A : in std_logic;  Y : out std_logic);

end IV_215;

architecture SYN_BEHAVIORAL of IV_215 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_214 is

   port( A : in std_logic;  Y : out std_logic);

end IV_214;

architecture SYN_BEHAVIORAL of IV_214 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_213 is

   port( A : in std_logic;  Y : out std_logic);

end IV_213;

architecture SYN_BEHAVIORAL of IV_213 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_212 is

   port( A : in std_logic;  Y : out std_logic);

end IV_212;

architecture SYN_BEHAVIORAL of IV_212 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_211 is

   port( A : in std_logic;  Y : out std_logic);

end IV_211;

architecture SYN_BEHAVIORAL of IV_211 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_210 is

   port( A : in std_logic;  Y : out std_logic);

end IV_210;

architecture SYN_BEHAVIORAL of IV_210 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_209 is

   port( A : in std_logic;  Y : out std_logic);

end IV_209;

architecture SYN_BEHAVIORAL of IV_209 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_208 is

   port( A : in std_logic;  Y : out std_logic);

end IV_208;

architecture SYN_BEHAVIORAL of IV_208 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_207 is

   port( A : in std_logic;  Y : out std_logic);

end IV_207;

architecture SYN_BEHAVIORAL of IV_207 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_206 is

   port( A : in std_logic;  Y : out std_logic);

end IV_206;

architecture SYN_BEHAVIORAL of IV_206 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_205 is

   port( A : in std_logic;  Y : out std_logic);

end IV_205;

architecture SYN_BEHAVIORAL of IV_205 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_204 is

   port( A : in std_logic;  Y : out std_logic);

end IV_204;

architecture SYN_BEHAVIORAL of IV_204 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_203 is

   port( A : in std_logic;  Y : out std_logic);

end IV_203;

architecture SYN_BEHAVIORAL of IV_203 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_202 is

   port( A : in std_logic;  Y : out std_logic);

end IV_202;

architecture SYN_BEHAVIORAL of IV_202 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_201 is

   port( A : in std_logic;  Y : out std_logic);

end IV_201;

architecture SYN_BEHAVIORAL of IV_201 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_200 is

   port( A : in std_logic;  Y : out std_logic);

end IV_200;

architecture SYN_BEHAVIORAL of IV_200 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_199 is

   port( A : in std_logic;  Y : out std_logic);

end IV_199;

architecture SYN_BEHAVIORAL of IV_199 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_198 is

   port( A : in std_logic;  Y : out std_logic);

end IV_198;

architecture SYN_BEHAVIORAL of IV_198 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_197 is

   port( A : in std_logic;  Y : out std_logic);

end IV_197;

architecture SYN_BEHAVIORAL of IV_197 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_196 is

   port( A : in std_logic;  Y : out std_logic);

end IV_196;

architecture SYN_BEHAVIORAL of IV_196 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_195 is

   port( A : in std_logic;  Y : out std_logic);

end IV_195;

architecture SYN_BEHAVIORAL of IV_195 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_194 is

   port( A : in std_logic;  Y : out std_logic);

end IV_194;

architecture SYN_BEHAVIORAL of IV_194 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_193 is

   port( A : in std_logic;  Y : out std_logic);

end IV_193;

architecture SYN_BEHAVIORAL of IV_193 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_192 is

   port( A : in std_logic;  Y : out std_logic);

end IV_192;

architecture SYN_BEHAVIORAL of IV_192 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_191 is

   port( A : in std_logic;  Y : out std_logic);

end IV_191;

architecture SYN_BEHAVIORAL of IV_191 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_190 is

   port( A : in std_logic;  Y : out std_logic);

end IV_190;

architecture SYN_BEHAVIORAL of IV_190 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_189 is

   port( A : in std_logic;  Y : out std_logic);

end IV_189;

architecture SYN_BEHAVIORAL of IV_189 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_188 is

   port( A : in std_logic;  Y : out std_logic);

end IV_188;

architecture SYN_BEHAVIORAL of IV_188 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_187 is

   port( A : in std_logic;  Y : out std_logic);

end IV_187;

architecture SYN_BEHAVIORAL of IV_187 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_186 is

   port( A : in std_logic;  Y : out std_logic);

end IV_186;

architecture SYN_BEHAVIORAL of IV_186 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_185 is

   port( A : in std_logic;  Y : out std_logic);

end IV_185;

architecture SYN_BEHAVIORAL of IV_185 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_184 is

   port( A : in std_logic;  Y : out std_logic);

end IV_184;

architecture SYN_BEHAVIORAL of IV_184 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_183 is

   port( A : in std_logic;  Y : out std_logic);

end IV_183;

architecture SYN_BEHAVIORAL of IV_183 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_182 is

   port( A : in std_logic;  Y : out std_logic);

end IV_182;

architecture SYN_BEHAVIORAL of IV_182 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_181 is

   port( A : in std_logic;  Y : out std_logic);

end IV_181;

architecture SYN_BEHAVIORAL of IV_181 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_180 is

   port( A : in std_logic;  Y : out std_logic);

end IV_180;

architecture SYN_BEHAVIORAL of IV_180 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_179 is

   port( A : in std_logic;  Y : out std_logic);

end IV_179;

architecture SYN_BEHAVIORAL of IV_179 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_178 is

   port( A : in std_logic;  Y : out std_logic);

end IV_178;

architecture SYN_BEHAVIORAL of IV_178 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_177 is

   port( A : in std_logic;  Y : out std_logic);

end IV_177;

architecture SYN_BEHAVIORAL of IV_177 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_176 is

   port( A : in std_logic;  Y : out std_logic);

end IV_176;

architecture SYN_BEHAVIORAL of IV_176 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_175 is

   port( A : in std_logic;  Y : out std_logic);

end IV_175;

architecture SYN_BEHAVIORAL of IV_175 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_174 is

   port( A : in std_logic;  Y : out std_logic);

end IV_174;

architecture SYN_BEHAVIORAL of IV_174 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_173 is

   port( A : in std_logic;  Y : out std_logic);

end IV_173;

architecture SYN_BEHAVIORAL of IV_173 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_172 is

   port( A : in std_logic;  Y : out std_logic);

end IV_172;

architecture SYN_BEHAVIORAL of IV_172 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_171 is

   port( A : in std_logic;  Y : out std_logic);

end IV_171;

architecture SYN_BEHAVIORAL of IV_171 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_170 is

   port( A : in std_logic;  Y : out std_logic);

end IV_170;

architecture SYN_BEHAVIORAL of IV_170 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_169 is

   port( A : in std_logic;  Y : out std_logic);

end IV_169;

architecture SYN_BEHAVIORAL of IV_169 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_168 is

   port( A : in std_logic;  Y : out std_logic);

end IV_168;

architecture SYN_BEHAVIORAL of IV_168 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_167 is

   port( A : in std_logic;  Y : out std_logic);

end IV_167;

architecture SYN_BEHAVIORAL of IV_167 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_166 is

   port( A : in std_logic;  Y : out std_logic);

end IV_166;

architecture SYN_BEHAVIORAL of IV_166 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_165 is

   port( A : in std_logic;  Y : out std_logic);

end IV_165;

architecture SYN_BEHAVIORAL of IV_165 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_164 is

   port( A : in std_logic;  Y : out std_logic);

end IV_164;

architecture SYN_BEHAVIORAL of IV_164 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_163 is

   port( A : in std_logic;  Y : out std_logic);

end IV_163;

architecture SYN_BEHAVIORAL of IV_163 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_162 is

   port( A : in std_logic;  Y : out std_logic);

end IV_162;

architecture SYN_BEHAVIORAL of IV_162 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_161 is

   port( A : in std_logic;  Y : out std_logic);

end IV_161;

architecture SYN_BEHAVIORAL of IV_161 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_160 is

   port( A : in std_logic;  Y : out std_logic);

end IV_160;

architecture SYN_BEHAVIORAL of IV_160 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_159 is

   port( A : in std_logic;  Y : out std_logic);

end IV_159;

architecture SYN_BEHAVIORAL of IV_159 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_158 is

   port( A : in std_logic;  Y : out std_logic);

end IV_158;

architecture SYN_BEHAVIORAL of IV_158 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_157 is

   port( A : in std_logic;  Y : out std_logic);

end IV_157;

architecture SYN_BEHAVIORAL of IV_157 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_156 is

   port( A : in std_logic;  Y : out std_logic);

end IV_156;

architecture SYN_BEHAVIORAL of IV_156 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_155 is

   port( A : in std_logic;  Y : out std_logic);

end IV_155;

architecture SYN_BEHAVIORAL of IV_155 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_154 is

   port( A : in std_logic;  Y : out std_logic);

end IV_154;

architecture SYN_BEHAVIORAL of IV_154 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_153 is

   port( A : in std_logic;  Y : out std_logic);

end IV_153;

architecture SYN_BEHAVIORAL of IV_153 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_152 is

   port( A : in std_logic;  Y : out std_logic);

end IV_152;

architecture SYN_BEHAVIORAL of IV_152 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_151 is

   port( A : in std_logic;  Y : out std_logic);

end IV_151;

architecture SYN_BEHAVIORAL of IV_151 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_150 is

   port( A : in std_logic;  Y : out std_logic);

end IV_150;

architecture SYN_BEHAVIORAL of IV_150 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_149 is

   port( A : in std_logic;  Y : out std_logic);

end IV_149;

architecture SYN_BEHAVIORAL of IV_149 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_148 is

   port( A : in std_logic;  Y : out std_logic);

end IV_148;

architecture SYN_BEHAVIORAL of IV_148 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_147 is

   port( A : in std_logic;  Y : out std_logic);

end IV_147;

architecture SYN_BEHAVIORAL of IV_147 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_146 is

   port( A : in std_logic;  Y : out std_logic);

end IV_146;

architecture SYN_BEHAVIORAL of IV_146 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_145 is

   port( A : in std_logic;  Y : out std_logic);

end IV_145;

architecture SYN_BEHAVIORAL of IV_145 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_144 is

   port( A : in std_logic;  Y : out std_logic);

end IV_144;

architecture SYN_BEHAVIORAL of IV_144 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_143 is

   port( A : in std_logic;  Y : out std_logic);

end IV_143;

architecture SYN_BEHAVIORAL of IV_143 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_142 is

   port( A : in std_logic;  Y : out std_logic);

end IV_142;

architecture SYN_BEHAVIORAL of IV_142 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_141 is

   port( A : in std_logic;  Y : out std_logic);

end IV_141;

architecture SYN_BEHAVIORAL of IV_141 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_140 is

   port( A : in std_logic;  Y : out std_logic);

end IV_140;

architecture SYN_BEHAVIORAL of IV_140 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_139 is

   port( A : in std_logic;  Y : out std_logic);

end IV_139;

architecture SYN_BEHAVIORAL of IV_139 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_138 is

   port( A : in std_logic;  Y : out std_logic);

end IV_138;

architecture SYN_BEHAVIORAL of IV_138 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_137 is

   port( A : in std_logic;  Y : out std_logic);

end IV_137;

architecture SYN_BEHAVIORAL of IV_137 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_136 is

   port( A : in std_logic;  Y : out std_logic);

end IV_136;

architecture SYN_BEHAVIORAL of IV_136 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_135 is

   port( A : in std_logic;  Y : out std_logic);

end IV_135;

architecture SYN_BEHAVIORAL of IV_135 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_134 is

   port( A : in std_logic;  Y : out std_logic);

end IV_134;

architecture SYN_BEHAVIORAL of IV_134 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_133 is

   port( A : in std_logic;  Y : out std_logic);

end IV_133;

architecture SYN_BEHAVIORAL of IV_133 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_132 is

   port( A : in std_logic;  Y : out std_logic);

end IV_132;

architecture SYN_BEHAVIORAL of IV_132 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_131 is

   port( A : in std_logic;  Y : out std_logic);

end IV_131;

architecture SYN_BEHAVIORAL of IV_131 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_130 is

   port( A : in std_logic;  Y : out std_logic);

end IV_130;

architecture SYN_BEHAVIORAL of IV_130 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_129 is

   port( A : in std_logic;  Y : out std_logic);

end IV_129;

architecture SYN_BEHAVIORAL of IV_129 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_128 is

   port( A : in std_logic;  Y : out std_logic);

end IV_128;

architecture SYN_BEHAVIORAL of IV_128 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_127 is

   port( A : in std_logic;  Y : out std_logic);

end IV_127;

architecture SYN_BEHAVIORAL of IV_127 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_126 is

   port( A : in std_logic;  Y : out std_logic);

end IV_126;

architecture SYN_BEHAVIORAL of IV_126 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_125 is

   port( A : in std_logic;  Y : out std_logic);

end IV_125;

architecture SYN_BEHAVIORAL of IV_125 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_124 is

   port( A : in std_logic;  Y : out std_logic);

end IV_124;

architecture SYN_BEHAVIORAL of IV_124 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_123 is

   port( A : in std_logic;  Y : out std_logic);

end IV_123;

architecture SYN_BEHAVIORAL of IV_123 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_122 is

   port( A : in std_logic;  Y : out std_logic);

end IV_122;

architecture SYN_BEHAVIORAL of IV_122 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_121 is

   port( A : in std_logic;  Y : out std_logic);

end IV_121;

architecture SYN_BEHAVIORAL of IV_121 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_120 is

   port( A : in std_logic;  Y : out std_logic);

end IV_120;

architecture SYN_BEHAVIORAL of IV_120 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_119 is

   port( A : in std_logic;  Y : out std_logic);

end IV_119;

architecture SYN_BEHAVIORAL of IV_119 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_118 is

   port( A : in std_logic;  Y : out std_logic);

end IV_118;

architecture SYN_BEHAVIORAL of IV_118 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_117 is

   port( A : in std_logic;  Y : out std_logic);

end IV_117;

architecture SYN_BEHAVIORAL of IV_117 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_116 is

   port( A : in std_logic;  Y : out std_logic);

end IV_116;

architecture SYN_BEHAVIORAL of IV_116 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_115 is

   port( A : in std_logic;  Y : out std_logic);

end IV_115;

architecture SYN_BEHAVIORAL of IV_115 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_114 is

   port( A : in std_logic;  Y : out std_logic);

end IV_114;

architecture SYN_BEHAVIORAL of IV_114 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_113 is

   port( A : in std_logic;  Y : out std_logic);

end IV_113;

architecture SYN_BEHAVIORAL of IV_113 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_112 is

   port( A : in std_logic;  Y : out std_logic);

end IV_112;

architecture SYN_BEHAVIORAL of IV_112 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_111 is

   port( A : in std_logic;  Y : out std_logic);

end IV_111;

architecture SYN_BEHAVIORAL of IV_111 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_110 is

   port( A : in std_logic;  Y : out std_logic);

end IV_110;

architecture SYN_BEHAVIORAL of IV_110 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_109 is

   port( A : in std_logic;  Y : out std_logic);

end IV_109;

architecture SYN_BEHAVIORAL of IV_109 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_108 is

   port( A : in std_logic;  Y : out std_logic);

end IV_108;

architecture SYN_BEHAVIORAL of IV_108 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_107 is

   port( A : in std_logic;  Y : out std_logic);

end IV_107;

architecture SYN_BEHAVIORAL of IV_107 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_106 is

   port( A : in std_logic;  Y : out std_logic);

end IV_106;

architecture SYN_BEHAVIORAL of IV_106 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_105 is

   port( A : in std_logic;  Y : out std_logic);

end IV_105;

architecture SYN_BEHAVIORAL of IV_105 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_104 is

   port( A : in std_logic;  Y : out std_logic);

end IV_104;

architecture SYN_BEHAVIORAL of IV_104 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_103 is

   port( A : in std_logic;  Y : out std_logic);

end IV_103;

architecture SYN_BEHAVIORAL of IV_103 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_102 is

   port( A : in std_logic;  Y : out std_logic);

end IV_102;

architecture SYN_BEHAVIORAL of IV_102 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_101 is

   port( A : in std_logic;  Y : out std_logic);

end IV_101;

architecture SYN_BEHAVIORAL of IV_101 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_100 is

   port( A : in std_logic;  Y : out std_logic);

end IV_100;

architecture SYN_BEHAVIORAL of IV_100 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_99 is

   port( A : in std_logic;  Y : out std_logic);

end IV_99;

architecture SYN_BEHAVIORAL of IV_99 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_98 is

   port( A : in std_logic;  Y : out std_logic);

end IV_98;

architecture SYN_BEHAVIORAL of IV_98 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_97 is

   port( A : in std_logic;  Y : out std_logic);

end IV_97;

architecture SYN_BEHAVIORAL of IV_97 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_96 is

   port( A : in std_logic;  Y : out std_logic);

end IV_96;

architecture SYN_BEHAVIORAL of IV_96 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_95 is

   port( A : in std_logic;  Y : out std_logic);

end IV_95;

architecture SYN_BEHAVIORAL of IV_95 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_94 is

   port( A : in std_logic;  Y : out std_logic);

end IV_94;

architecture SYN_BEHAVIORAL of IV_94 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_93 is

   port( A : in std_logic;  Y : out std_logic);

end IV_93;

architecture SYN_BEHAVIORAL of IV_93 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_92 is

   port( A : in std_logic;  Y : out std_logic);

end IV_92;

architecture SYN_BEHAVIORAL of IV_92 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_91 is

   port( A : in std_logic;  Y : out std_logic);

end IV_91;

architecture SYN_BEHAVIORAL of IV_91 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_90 is

   port( A : in std_logic;  Y : out std_logic);

end IV_90;

architecture SYN_BEHAVIORAL of IV_90 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_89 is

   port( A : in std_logic;  Y : out std_logic);

end IV_89;

architecture SYN_BEHAVIORAL of IV_89 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_88 is

   port( A : in std_logic;  Y : out std_logic);

end IV_88;

architecture SYN_BEHAVIORAL of IV_88 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_87 is

   port( A : in std_logic;  Y : out std_logic);

end IV_87;

architecture SYN_BEHAVIORAL of IV_87 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_86 is

   port( A : in std_logic;  Y : out std_logic);

end IV_86;

architecture SYN_BEHAVIORAL of IV_86 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_85 is

   port( A : in std_logic;  Y : out std_logic);

end IV_85;

architecture SYN_BEHAVIORAL of IV_85 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_84 is

   port( A : in std_logic;  Y : out std_logic);

end IV_84;

architecture SYN_BEHAVIORAL of IV_84 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_83 is

   port( A : in std_logic;  Y : out std_logic);

end IV_83;

architecture SYN_BEHAVIORAL of IV_83 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_82 is

   port( A : in std_logic;  Y : out std_logic);

end IV_82;

architecture SYN_BEHAVIORAL of IV_82 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_81 is

   port( A : in std_logic;  Y : out std_logic);

end IV_81;

architecture SYN_BEHAVIORAL of IV_81 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_80 is

   port( A : in std_logic;  Y : out std_logic);

end IV_80;

architecture SYN_BEHAVIORAL of IV_80 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_79 is

   port( A : in std_logic;  Y : out std_logic);

end IV_79;

architecture SYN_BEHAVIORAL of IV_79 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_78 is

   port( A : in std_logic;  Y : out std_logic);

end IV_78;

architecture SYN_BEHAVIORAL of IV_78 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_77 is

   port( A : in std_logic;  Y : out std_logic);

end IV_77;

architecture SYN_BEHAVIORAL of IV_77 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_76 is

   port( A : in std_logic;  Y : out std_logic);

end IV_76;

architecture SYN_BEHAVIORAL of IV_76 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_75 is

   port( A : in std_logic;  Y : out std_logic);

end IV_75;

architecture SYN_BEHAVIORAL of IV_75 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_74 is

   port( A : in std_logic;  Y : out std_logic);

end IV_74;

architecture SYN_BEHAVIORAL of IV_74 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_73 is

   port( A : in std_logic;  Y : out std_logic);

end IV_73;

architecture SYN_BEHAVIORAL of IV_73 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_72 is

   port( A : in std_logic;  Y : out std_logic);

end IV_72;

architecture SYN_BEHAVIORAL of IV_72 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_71 is

   port( A : in std_logic;  Y : out std_logic);

end IV_71;

architecture SYN_BEHAVIORAL of IV_71 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_70 is

   port( A : in std_logic;  Y : out std_logic);

end IV_70;

architecture SYN_BEHAVIORAL of IV_70 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_69 is

   port( A : in std_logic;  Y : out std_logic);

end IV_69;

architecture SYN_BEHAVIORAL of IV_69 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_68 is

   port( A : in std_logic;  Y : out std_logic);

end IV_68;

architecture SYN_BEHAVIORAL of IV_68 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_67 is

   port( A : in std_logic;  Y : out std_logic);

end IV_67;

architecture SYN_BEHAVIORAL of IV_67 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_66 is

   port( A : in std_logic;  Y : out std_logic);

end IV_66;

architecture SYN_BEHAVIORAL of IV_66 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_65 is

   port( A : in std_logic;  Y : out std_logic);

end IV_65;

architecture SYN_BEHAVIORAL of IV_65 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_64 is

   port( A : in std_logic;  Y : out std_logic);

end IV_64;

architecture SYN_BEHAVIORAL of IV_64 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_63 is

   port( A : in std_logic;  Y : out std_logic);

end IV_63;

architecture SYN_BEHAVIORAL of IV_63 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_62 is

   port( A : in std_logic;  Y : out std_logic);

end IV_62;

architecture SYN_BEHAVIORAL of IV_62 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_61 is

   port( A : in std_logic;  Y : out std_logic);

end IV_61;

architecture SYN_BEHAVIORAL of IV_61 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_60 is

   port( A : in std_logic;  Y : out std_logic);

end IV_60;

architecture SYN_BEHAVIORAL of IV_60 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_59 is

   port( A : in std_logic;  Y : out std_logic);

end IV_59;

architecture SYN_BEHAVIORAL of IV_59 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_58 is

   port( A : in std_logic;  Y : out std_logic);

end IV_58;

architecture SYN_BEHAVIORAL of IV_58 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_57 is

   port( A : in std_logic;  Y : out std_logic);

end IV_57;

architecture SYN_BEHAVIORAL of IV_57 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_56 is

   port( A : in std_logic;  Y : out std_logic);

end IV_56;

architecture SYN_BEHAVIORAL of IV_56 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_55 is

   port( A : in std_logic;  Y : out std_logic);

end IV_55;

architecture SYN_BEHAVIORAL of IV_55 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_54 is

   port( A : in std_logic;  Y : out std_logic);

end IV_54;

architecture SYN_BEHAVIORAL of IV_54 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_53 is

   port( A : in std_logic;  Y : out std_logic);

end IV_53;

architecture SYN_BEHAVIORAL of IV_53 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_52 is

   port( A : in std_logic;  Y : out std_logic);

end IV_52;

architecture SYN_BEHAVIORAL of IV_52 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_51 is

   port( A : in std_logic;  Y : out std_logic);

end IV_51;

architecture SYN_BEHAVIORAL of IV_51 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_50 is

   port( A : in std_logic;  Y : out std_logic);

end IV_50;

architecture SYN_BEHAVIORAL of IV_50 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_49 is

   port( A : in std_logic;  Y : out std_logic);

end IV_49;

architecture SYN_BEHAVIORAL of IV_49 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_48 is

   port( A : in std_logic;  Y : out std_logic);

end IV_48;

architecture SYN_BEHAVIORAL of IV_48 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_47 is

   port( A : in std_logic;  Y : out std_logic);

end IV_47;

architecture SYN_BEHAVIORAL of IV_47 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_46 is

   port( A : in std_logic;  Y : out std_logic);

end IV_46;

architecture SYN_BEHAVIORAL of IV_46 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_45 is

   port( A : in std_logic;  Y : out std_logic);

end IV_45;

architecture SYN_BEHAVIORAL of IV_45 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_44 is

   port( A : in std_logic;  Y : out std_logic);

end IV_44;

architecture SYN_BEHAVIORAL of IV_44 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_43 is

   port( A : in std_logic;  Y : out std_logic);

end IV_43;

architecture SYN_BEHAVIORAL of IV_43 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_42 is

   port( A : in std_logic;  Y : out std_logic);

end IV_42;

architecture SYN_BEHAVIORAL of IV_42 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_41 is

   port( A : in std_logic;  Y : out std_logic);

end IV_41;

architecture SYN_BEHAVIORAL of IV_41 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_40 is

   port( A : in std_logic;  Y : out std_logic);

end IV_40;

architecture SYN_BEHAVIORAL of IV_40 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_39 is

   port( A : in std_logic;  Y : out std_logic);

end IV_39;

architecture SYN_BEHAVIORAL of IV_39 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_38 is

   port( A : in std_logic;  Y : out std_logic);

end IV_38;

architecture SYN_BEHAVIORAL of IV_38 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_37 is

   port( A : in std_logic;  Y : out std_logic);

end IV_37;

architecture SYN_BEHAVIORAL of IV_37 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_36 is

   port( A : in std_logic;  Y : out std_logic);

end IV_36;

architecture SYN_BEHAVIORAL of IV_36 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_35 is

   port( A : in std_logic;  Y : out std_logic);

end IV_35;

architecture SYN_BEHAVIORAL of IV_35 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_34 is

   port( A : in std_logic;  Y : out std_logic);

end IV_34;

architecture SYN_BEHAVIORAL of IV_34 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_33 is

   port( A : in std_logic;  Y : out std_logic);

end IV_33;

architecture SYN_BEHAVIORAL of IV_33 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_32 is

   port( A : in std_logic;  Y : out std_logic);

end IV_32;

architecture SYN_BEHAVIORAL of IV_32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_31 is

   port( A : in std_logic;  Y : out std_logic);

end IV_31;

architecture SYN_BEHAVIORAL of IV_31 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_30 is

   port( A : in std_logic;  Y : out std_logic);

end IV_30;

architecture SYN_BEHAVIORAL of IV_30 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_29 is

   port( A : in std_logic;  Y : out std_logic);

end IV_29;

architecture SYN_BEHAVIORAL of IV_29 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_28 is

   port( A : in std_logic;  Y : out std_logic);

end IV_28;

architecture SYN_BEHAVIORAL of IV_28 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_27 is

   port( A : in std_logic;  Y : out std_logic);

end IV_27;

architecture SYN_BEHAVIORAL of IV_27 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_26 is

   port( A : in std_logic;  Y : out std_logic);

end IV_26;

architecture SYN_BEHAVIORAL of IV_26 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_25 is

   port( A : in std_logic;  Y : out std_logic);

end IV_25;

architecture SYN_BEHAVIORAL of IV_25 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_24 is

   port( A : in std_logic;  Y : out std_logic);

end IV_24;

architecture SYN_BEHAVIORAL of IV_24 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_23 is

   port( A : in std_logic;  Y : out std_logic);

end IV_23;

architecture SYN_BEHAVIORAL of IV_23 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_22 is

   port( A : in std_logic;  Y : out std_logic);

end IV_22;

architecture SYN_BEHAVIORAL of IV_22 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_21 is

   port( A : in std_logic;  Y : out std_logic);

end IV_21;

architecture SYN_BEHAVIORAL of IV_21 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_20 is

   port( A : in std_logic;  Y : out std_logic);

end IV_20;

architecture SYN_BEHAVIORAL of IV_20 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_19 is

   port( A : in std_logic;  Y : out std_logic);

end IV_19;

architecture SYN_BEHAVIORAL of IV_19 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_18 is

   port( A : in std_logic;  Y : out std_logic);

end IV_18;

architecture SYN_BEHAVIORAL of IV_18 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_17 is

   port( A : in std_logic;  Y : out std_logic);

end IV_17;

architecture SYN_BEHAVIORAL of IV_17 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_16 is

   port( A : in std_logic;  Y : out std_logic);

end IV_16;

architecture SYN_BEHAVIORAL of IV_16 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_15 is

   port( A : in std_logic;  Y : out std_logic);

end IV_15;

architecture SYN_BEHAVIORAL of IV_15 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_14 is

   port( A : in std_logic;  Y : out std_logic);

end IV_14;

architecture SYN_BEHAVIORAL of IV_14 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_13 is

   port( A : in std_logic;  Y : out std_logic);

end IV_13;

architecture SYN_BEHAVIORAL of IV_13 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_12 is

   port( A : in std_logic;  Y : out std_logic);

end IV_12;

architecture SYN_BEHAVIORAL of IV_12 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_11 is

   port( A : in std_logic;  Y : out std_logic);

end IV_11;

architecture SYN_BEHAVIORAL of IV_11 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_10 is

   port( A : in std_logic;  Y : out std_logic);

end IV_10;

architecture SYN_BEHAVIORAL of IV_10 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_9 is

   port( A : in std_logic;  Y : out std_logic);

end IV_9;

architecture SYN_BEHAVIORAL of IV_9 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_8 is

   port( A : in std_logic;  Y : out std_logic);

end IV_8;

architecture SYN_BEHAVIORAL of IV_8 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_7 is

   port( A : in std_logic;  Y : out std_logic);

end IV_7;

architecture SYN_BEHAVIORAL of IV_7 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_6 is

   port( A : in std_logic;  Y : out std_logic);

end IV_6;

architecture SYN_BEHAVIORAL of IV_6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_5 is

   port( A : in std_logic;  Y : out std_logic);

end IV_5;

architecture SYN_BEHAVIORAL of IV_5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_4 is

   port( A : in std_logic;  Y : out std_logic);

end IV_4;

architecture SYN_BEHAVIORAL of IV_4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_3 is

   port( A : in std_logic;  Y : out std_logic);

end IV_3;

architecture SYN_BEHAVIORAL of IV_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_2 is

   port( A : in std_logic;  Y : out std_logic);

end IV_2;

architecture SYN_BEHAVIORAL of IV_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_1 is

   port( A : in std_logic;  Y : out std_logic);

end IV_1;

architecture SYN_BEHAVIORAL of IV_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_255 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_255;

architecture SYN_STRUCTURAL of MUX21_255 is

   component ND2_763
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_764
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_765
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_255
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_255 port map( A => S, Y => SB);
   UND1 : ND2_765 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_764 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_763 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_254 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_254;

architecture SYN_STRUCTURAL of MUX21_254 is

   component ND2_760
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_761
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_762
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_254
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_254 port map( A => S, Y => SB);
   UND1 : ND2_762 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_761 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_760 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_253 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_253;

architecture SYN_STRUCTURAL of MUX21_253 is

   component ND2_757
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_758
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_759
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_253
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_253 port map( A => S, Y => SB);
   UND1 : ND2_759 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_758 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_757 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_252 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_252;

architecture SYN_STRUCTURAL of MUX21_252 is

   component ND2_754
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_755
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_756
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_252
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_252 port map( A => S, Y => SB);
   UND1 : ND2_756 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_755 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_754 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_251 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_251;

architecture SYN_STRUCTURAL of MUX21_251 is

   component ND2_751
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_752
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_753
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_251
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_251 port map( A => S, Y => SB);
   UND1 : ND2_753 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_752 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_751 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_250 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_250;

architecture SYN_STRUCTURAL of MUX21_250 is

   component ND2_748
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_749
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_750
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_250
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_250 port map( A => S, Y => SB);
   UND1 : ND2_750 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_749 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_748 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_249 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_249;

architecture SYN_STRUCTURAL of MUX21_249 is

   component ND2_745
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_746
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_747
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_249
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_249 port map( A => S, Y => SB);
   UND1 : ND2_747 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_746 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_745 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_248 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_248;

architecture SYN_STRUCTURAL of MUX21_248 is

   component ND2_742
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_743
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_744
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_248
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_248 port map( A => S, Y => SB);
   UND1 : ND2_744 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_743 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_742 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_247 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_247;

architecture SYN_STRUCTURAL of MUX21_247 is

   component ND2_739
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_740
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_741
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_247
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_247 port map( A => S, Y => SB);
   UND1 : ND2_741 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_740 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_739 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_246 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_246;

architecture SYN_STRUCTURAL of MUX21_246 is

   component ND2_736
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_737
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_738
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_246
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_246 port map( A => S, Y => SB);
   UND1 : ND2_738 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_737 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_736 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_245 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_245;

architecture SYN_STRUCTURAL of MUX21_245 is

   component ND2_733
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_734
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_735
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_245
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_245 port map( A => S, Y => SB);
   UND1 : ND2_735 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_734 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_733 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_244 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_244;

architecture SYN_STRUCTURAL of MUX21_244 is

   component ND2_730
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_731
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_732
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_244
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_244 port map( A => S, Y => SB);
   UND1 : ND2_732 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_731 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_730 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_243 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_243;

architecture SYN_STRUCTURAL of MUX21_243 is

   component ND2_727
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_728
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_729
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_243
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_243 port map( A => S, Y => SB);
   UND1 : ND2_729 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_728 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_727 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_242 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_242;

architecture SYN_STRUCTURAL of MUX21_242 is

   component ND2_724
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_725
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_726
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_242
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_242 port map( A => S, Y => SB);
   UND1 : ND2_726 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_725 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_724 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_241 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_241;

architecture SYN_STRUCTURAL of MUX21_241 is

   component ND2_721
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_722
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_723
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_241
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_241 port map( A => S, Y => SB);
   UND1 : ND2_723 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_722 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_721 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_240 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_240;

architecture SYN_STRUCTURAL of MUX21_240 is

   component ND2_718
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_719
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_720
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_240
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_240 port map( A => S, Y => SB);
   UND1 : ND2_720 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_719 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_718 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_239 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_239;

architecture SYN_STRUCTURAL of MUX21_239 is

   component ND2_715
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_716
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_717
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_239
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_239 port map( A => S, Y => SB);
   UND1 : ND2_717 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_716 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_715 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_238 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_238;

architecture SYN_STRUCTURAL of MUX21_238 is

   component ND2_712
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_713
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_714
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_238
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_238 port map( A => S, Y => SB);
   UND1 : ND2_714 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_713 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_712 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_237 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_237;

architecture SYN_STRUCTURAL of MUX21_237 is

   component ND2_709
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_710
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_711
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_237
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_237 port map( A => S, Y => SB);
   UND1 : ND2_711 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_710 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_709 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_236 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_236;

architecture SYN_STRUCTURAL of MUX21_236 is

   component ND2_706
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_707
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_708
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_236
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_236 port map( A => S, Y => SB);
   UND1 : ND2_708 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_707 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_706 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_235 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_235;

architecture SYN_STRUCTURAL of MUX21_235 is

   component ND2_703
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_704
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_705
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_235
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_235 port map( A => S, Y => SB);
   UND1 : ND2_705 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_704 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_703 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_234 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_234;

architecture SYN_STRUCTURAL of MUX21_234 is

   component ND2_700
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_701
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_702
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_234
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_234 port map( A => S, Y => SB);
   UND1 : ND2_702 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_701 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_700 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_233 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_233;

architecture SYN_STRUCTURAL of MUX21_233 is

   component ND2_697
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_698
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_699
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_233
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_233 port map( A => S, Y => SB);
   UND1 : ND2_699 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_698 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_697 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_232 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_232;

architecture SYN_STRUCTURAL of MUX21_232 is

   component ND2_694
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_695
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_696
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_232
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_232 port map( A => S, Y => SB);
   UND1 : ND2_696 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_695 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_694 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_231 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_231;

architecture SYN_STRUCTURAL of MUX21_231 is

   component ND2_691
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_692
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_693
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_231
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_231 port map( A => S, Y => SB);
   UND1 : ND2_693 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_692 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_691 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_230 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_230;

architecture SYN_STRUCTURAL of MUX21_230 is

   component ND2_688
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_689
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_690
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_230
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_230 port map( A => S, Y => SB);
   UND1 : ND2_690 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_689 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_688 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_229 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_229;

architecture SYN_STRUCTURAL of MUX21_229 is

   component ND2_685
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_686
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_687
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_229
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_229 port map( A => S, Y => SB);
   UND1 : ND2_687 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_686 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_685 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_228 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_228;

architecture SYN_STRUCTURAL of MUX21_228 is

   component ND2_682
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_683
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_684
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_228
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_228 port map( A => S, Y => SB);
   UND1 : ND2_684 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_683 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_682 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_227 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_227;

architecture SYN_STRUCTURAL of MUX21_227 is

   component ND2_679
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_680
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_681
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_227
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_227 port map( A => S, Y => SB);
   UND1 : ND2_681 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_680 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_679 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_226 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_226;

architecture SYN_STRUCTURAL of MUX21_226 is

   component ND2_676
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_677
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_678
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_226
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_226 port map( A => S, Y => SB);
   UND1 : ND2_678 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_677 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_676 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_225 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_225;

architecture SYN_STRUCTURAL of MUX21_225 is

   component ND2_673
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_674
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_675
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_225
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_225 port map( A => S, Y => SB);
   UND1 : ND2_675 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_674 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_673 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_224 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_224;

architecture SYN_STRUCTURAL of MUX21_224 is

   component ND2_670
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_671
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_672
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_224
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_224 port map( A => S, Y => SB);
   UND1 : ND2_672 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_671 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_670 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_223 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_223;

architecture SYN_STRUCTURAL of MUX21_223 is

   component ND2_667
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_668
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_669
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_223
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_223 port map( A => S, Y => SB);
   UND1 : ND2_669 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_668 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_667 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_222 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_222;

architecture SYN_STRUCTURAL of MUX21_222 is

   component ND2_664
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_665
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_666
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_222
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_222 port map( A => S, Y => SB);
   UND1 : ND2_666 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_665 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_664 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_221 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_221;

architecture SYN_STRUCTURAL of MUX21_221 is

   component ND2_661
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_662
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_663
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_221
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_221 port map( A => S, Y => SB);
   UND1 : ND2_663 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_662 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_661 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_220 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_220;

architecture SYN_STRUCTURAL of MUX21_220 is

   component ND2_658
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_659
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_660
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_220
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_220 port map( A => S, Y => SB);
   UND1 : ND2_660 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_659 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_658 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_219 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_219;

architecture SYN_STRUCTURAL of MUX21_219 is

   component ND2_655
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_656
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_657
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_219
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_219 port map( A => S, Y => SB);
   UND1 : ND2_657 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_656 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_655 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_218 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_218;

architecture SYN_STRUCTURAL of MUX21_218 is

   component ND2_652
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_653
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_654
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_218
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_218 port map( A => S, Y => SB);
   UND1 : ND2_654 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_653 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_652 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_217 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_217;

architecture SYN_STRUCTURAL of MUX21_217 is

   component ND2_649
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_650
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_651
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_217
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_217 port map( A => S, Y => SB);
   UND1 : ND2_651 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_650 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_649 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_216 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_216;

architecture SYN_STRUCTURAL of MUX21_216 is

   component ND2_646
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_647
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_648
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_216
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_216 port map( A => S, Y => SB);
   UND1 : ND2_648 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_647 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_646 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_215 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_215;

architecture SYN_STRUCTURAL of MUX21_215 is

   component ND2_643
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_644
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_645
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_215
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_215 port map( A => S, Y => SB);
   UND1 : ND2_645 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_644 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_643 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_214 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_214;

architecture SYN_STRUCTURAL of MUX21_214 is

   component ND2_640
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_641
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_642
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_214
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_214 port map( A => S, Y => SB);
   UND1 : ND2_642 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_641 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_640 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_213 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_213;

architecture SYN_STRUCTURAL of MUX21_213 is

   component ND2_637
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_638
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_639
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_213
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_213 port map( A => S, Y => SB);
   UND1 : ND2_639 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_638 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_637 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_212 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_212;

architecture SYN_STRUCTURAL of MUX21_212 is

   component ND2_634
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_635
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_636
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_212
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_212 port map( A => S, Y => SB);
   UND1 : ND2_636 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_635 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_634 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_211 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_211;

architecture SYN_STRUCTURAL of MUX21_211 is

   component ND2_631
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_632
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_633
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_211
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_211 port map( A => S, Y => SB);
   UND1 : ND2_633 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_632 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_631 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_210 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_210;

architecture SYN_STRUCTURAL of MUX21_210 is

   component ND2_628
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_629
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_630
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_210
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_210 port map( A => S, Y => SB);
   UND1 : ND2_630 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_629 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_628 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_209 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_209;

architecture SYN_STRUCTURAL of MUX21_209 is

   component ND2_625
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_626
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_627
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_209
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_209 port map( A => S, Y => SB);
   UND1 : ND2_627 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_626 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_625 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_208 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_208;

architecture SYN_STRUCTURAL of MUX21_208 is

   component ND2_622
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_623
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_624
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_208
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_208 port map( A => S, Y => SB);
   UND1 : ND2_624 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_623 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_622 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_207 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_207;

architecture SYN_STRUCTURAL of MUX21_207 is

   component ND2_619
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_620
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_621
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_207
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_207 port map( A => S, Y => SB);
   UND1 : ND2_621 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_620 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_619 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_206 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_206;

architecture SYN_STRUCTURAL of MUX21_206 is

   component ND2_616
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_617
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_618
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_206
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_206 port map( A => S, Y => SB);
   UND1 : ND2_618 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_617 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_616 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_205 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_205;

architecture SYN_STRUCTURAL of MUX21_205 is

   component ND2_613
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_614
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_615
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_205
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_205 port map( A => S, Y => SB);
   UND1 : ND2_615 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_614 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_613 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_204 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_204;

architecture SYN_STRUCTURAL of MUX21_204 is

   component ND2_610
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_611
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_612
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_204
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_204 port map( A => S, Y => SB);
   UND1 : ND2_612 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_611 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_610 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_203 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_203;

architecture SYN_STRUCTURAL of MUX21_203 is

   component ND2_607
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_608
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_609
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_203
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_203 port map( A => S, Y => SB);
   UND1 : ND2_609 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_608 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_607 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_202 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_202;

architecture SYN_STRUCTURAL of MUX21_202 is

   component ND2_604
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_605
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_606
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_202
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_202 port map( A => S, Y => SB);
   UND1 : ND2_606 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_605 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_604 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_201 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_201;

architecture SYN_STRUCTURAL of MUX21_201 is

   component ND2_601
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_602
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_603
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_201
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_201 port map( A => S, Y => SB);
   UND1 : ND2_603 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_602 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_601 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_200 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_200;

architecture SYN_STRUCTURAL of MUX21_200 is

   component ND2_598
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_599
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_600
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_200
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_200 port map( A => S, Y => SB);
   UND1 : ND2_600 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_599 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_598 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_199 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_199;

architecture SYN_STRUCTURAL of MUX21_199 is

   component ND2_595
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_596
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_597
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_199
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_199 port map( A => S, Y => SB);
   UND1 : ND2_597 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_596 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_595 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_198 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_198;

architecture SYN_STRUCTURAL of MUX21_198 is

   component ND2_592
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_593
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_594
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_198
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_198 port map( A => S, Y => SB);
   UND1 : ND2_594 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_593 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_592 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_197 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_197;

architecture SYN_STRUCTURAL of MUX21_197 is

   component ND2_589
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_590
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_591
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_197
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_197 port map( A => S, Y => SB);
   UND1 : ND2_591 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_590 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_589 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_196 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_196;

architecture SYN_STRUCTURAL of MUX21_196 is

   component ND2_586
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_587
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_588
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_196
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_196 port map( A => S, Y => SB);
   UND1 : ND2_588 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_587 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_586 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_195 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_195;

architecture SYN_STRUCTURAL of MUX21_195 is

   component ND2_583
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_584
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_585
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_195
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_195 port map( A => S, Y => SB);
   UND1 : ND2_585 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_584 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_583 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_194 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_194;

architecture SYN_STRUCTURAL of MUX21_194 is

   component ND2_580
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_581
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_582
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_194
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_194 port map( A => S, Y => SB);
   UND1 : ND2_582 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_581 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_580 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_193 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_193;

architecture SYN_STRUCTURAL of MUX21_193 is

   component ND2_577
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_578
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_579
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_193
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_193 port map( A => S, Y => SB);
   UND1 : ND2_579 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_578 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_577 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_192 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_192;

architecture SYN_STRUCTURAL of MUX21_192 is

   component ND2_574
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_575
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_576
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_192
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_192 port map( A => S, Y => SB);
   UND1 : ND2_576 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_575 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_574 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_191 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_191;

architecture SYN_STRUCTURAL of MUX21_191 is

   component ND2_571
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_572
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_573
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_191
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_191 port map( A => S, Y => SB);
   UND1 : ND2_573 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_572 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_571 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_190 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_190;

architecture SYN_STRUCTURAL of MUX21_190 is

   component ND2_568
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_569
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_570
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_190
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_190 port map( A => S, Y => SB);
   UND1 : ND2_570 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_569 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_568 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_189 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_189;

architecture SYN_STRUCTURAL of MUX21_189 is

   component ND2_565
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_566
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_567
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_189
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_189 port map( A => S, Y => SB);
   UND1 : ND2_567 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_566 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_565 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_188 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_188;

architecture SYN_STRUCTURAL of MUX21_188 is

   component ND2_562
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_563
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_564
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_188
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_188 port map( A => S, Y => SB);
   UND1 : ND2_564 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_563 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_562 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_187 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_187;

architecture SYN_STRUCTURAL of MUX21_187 is

   component ND2_559
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_560
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_561
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_187
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_187 port map( A => S, Y => SB);
   UND1 : ND2_561 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_560 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_559 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_186 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_186;

architecture SYN_STRUCTURAL of MUX21_186 is

   component ND2_556
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_557
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_558
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_186
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_186 port map( A => S, Y => SB);
   UND1 : ND2_558 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_557 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_556 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_185 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_185;

architecture SYN_STRUCTURAL of MUX21_185 is

   component ND2_553
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_554
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_555
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_185
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_185 port map( A => S, Y => SB);
   UND1 : ND2_555 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_554 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_553 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_184 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_184;

architecture SYN_STRUCTURAL of MUX21_184 is

   component ND2_550
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_551
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_552
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_184
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_184 port map( A => S, Y => SB);
   UND1 : ND2_552 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_551 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_550 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_183 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_183;

architecture SYN_STRUCTURAL of MUX21_183 is

   component ND2_547
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_548
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_549
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_183
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_183 port map( A => S, Y => SB);
   UND1 : ND2_549 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_548 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_547 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_182 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_182;

architecture SYN_STRUCTURAL of MUX21_182 is

   component ND2_544
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_545
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_546
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_182
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_182 port map( A => S, Y => SB);
   UND1 : ND2_546 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_545 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_544 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_181 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_181;

architecture SYN_STRUCTURAL of MUX21_181 is

   component ND2_541
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_542
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_543
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_181
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_181 port map( A => S, Y => SB);
   UND1 : ND2_543 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_542 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_541 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_180 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_180;

architecture SYN_STRUCTURAL of MUX21_180 is

   component ND2_538
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_539
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_540
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_180
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_180 port map( A => S, Y => SB);
   UND1 : ND2_540 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_539 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_538 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_179 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_179;

architecture SYN_STRUCTURAL of MUX21_179 is

   component ND2_535
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_536
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_537
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_179
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_179 port map( A => S, Y => SB);
   UND1 : ND2_537 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_536 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_535 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_178 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_178;

architecture SYN_STRUCTURAL of MUX21_178 is

   component ND2_532
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_533
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_534
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_178
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_178 port map( A => S, Y => SB);
   UND1 : ND2_534 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_533 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_532 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_177 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_177;

architecture SYN_STRUCTURAL of MUX21_177 is

   component ND2_529
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_530
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_531
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_177
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_177 port map( A => S, Y => SB);
   UND1 : ND2_531 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_530 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_529 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_176 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_176;

architecture SYN_STRUCTURAL of MUX21_176 is

   component ND2_526
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_527
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_528
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_176
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_176 port map( A => S, Y => SB);
   UND1 : ND2_528 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_527 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_526 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_175 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_175;

architecture SYN_STRUCTURAL of MUX21_175 is

   component ND2_523
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_524
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_525
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_175
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_175 port map( A => S, Y => SB);
   UND1 : ND2_525 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_524 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_523 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_174 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_174;

architecture SYN_STRUCTURAL of MUX21_174 is

   component ND2_520
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_521
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_522
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_174
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_174 port map( A => S, Y => SB);
   UND1 : ND2_522 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_521 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_520 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_173 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_173;

architecture SYN_STRUCTURAL of MUX21_173 is

   component ND2_517
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_518
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_519
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_173
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_173 port map( A => S, Y => SB);
   UND1 : ND2_519 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_518 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_517 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_172 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_172;

architecture SYN_STRUCTURAL of MUX21_172 is

   component ND2_514
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_515
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_516
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_172
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_172 port map( A => S, Y => SB);
   UND1 : ND2_516 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_515 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_514 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_171 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_171;

architecture SYN_STRUCTURAL of MUX21_171 is

   component ND2_511
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_512
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_513
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_171
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_171 port map( A => S, Y => SB);
   UND1 : ND2_513 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_512 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_511 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_170 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_170;

architecture SYN_STRUCTURAL of MUX21_170 is

   component ND2_508
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_509
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_510
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_170
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_170 port map( A => S, Y => SB);
   UND1 : ND2_510 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_509 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_508 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_169 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_169;

architecture SYN_STRUCTURAL of MUX21_169 is

   component ND2_505
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_506
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_507
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_169
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_169 port map( A => S, Y => SB);
   UND1 : ND2_507 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_506 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_505 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_168 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_168;

architecture SYN_STRUCTURAL of MUX21_168 is

   component ND2_502
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_503
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_504
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_168
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_168 port map( A => S, Y => SB);
   UND1 : ND2_504 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_503 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_502 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_167 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_167;

architecture SYN_STRUCTURAL of MUX21_167 is

   component ND2_499
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_500
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_501
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_167
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_167 port map( A => S, Y => SB);
   UND1 : ND2_501 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_500 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_499 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_166 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_166;

architecture SYN_STRUCTURAL of MUX21_166 is

   component ND2_496
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_497
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_498
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_166
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_166 port map( A => S, Y => SB);
   UND1 : ND2_498 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_497 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_496 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_165 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_165;

architecture SYN_STRUCTURAL of MUX21_165 is

   component ND2_493
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_494
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_495
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_165
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_165 port map( A => S, Y => SB);
   UND1 : ND2_495 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_494 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_493 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_164 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_164;

architecture SYN_STRUCTURAL of MUX21_164 is

   component ND2_490
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_491
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_492
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_164
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_164 port map( A => S, Y => SB);
   UND1 : ND2_492 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_491 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_490 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_163 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_163;

architecture SYN_STRUCTURAL of MUX21_163 is

   component ND2_487
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_488
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_489
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_163
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_163 port map( A => S, Y => SB);
   UND1 : ND2_489 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_488 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_487 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_162 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_162;

architecture SYN_STRUCTURAL of MUX21_162 is

   component ND2_484
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_485
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_486
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_162
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_162 port map( A => S, Y => SB);
   UND1 : ND2_486 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_485 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_484 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_161 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_161;

architecture SYN_STRUCTURAL of MUX21_161 is

   component ND2_481
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_482
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_483
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_161
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_161 port map( A => S, Y => SB);
   UND1 : ND2_483 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_482 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_481 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_160 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_160;

architecture SYN_STRUCTURAL of MUX21_160 is

   component ND2_478
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_479
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_480
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_160
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_160 port map( A => S, Y => SB);
   UND1 : ND2_480 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_479 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_478 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_159 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_159;

architecture SYN_STRUCTURAL of MUX21_159 is

   component ND2_475
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_476
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_477
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_159
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_159 port map( A => S, Y => SB);
   UND1 : ND2_477 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_476 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_475 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_158 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_158;

architecture SYN_STRUCTURAL of MUX21_158 is

   component ND2_472
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_473
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_474
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_158
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_158 port map( A => S, Y => SB);
   UND1 : ND2_474 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_473 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_472 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_157 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_157;

architecture SYN_STRUCTURAL of MUX21_157 is

   component ND2_469
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_470
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_471
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_157
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_157 port map( A => S, Y => SB);
   UND1 : ND2_471 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_470 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_469 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_156 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_156;

architecture SYN_STRUCTURAL of MUX21_156 is

   component ND2_466
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_467
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_468
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_156
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_156 port map( A => S, Y => SB);
   UND1 : ND2_468 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_467 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_466 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_155 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_155;

architecture SYN_STRUCTURAL of MUX21_155 is

   component ND2_463
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_464
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_465
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_155
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_155 port map( A => S, Y => SB);
   UND1 : ND2_465 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_464 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_463 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_154 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_154;

architecture SYN_STRUCTURAL of MUX21_154 is

   component ND2_460
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_461
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_462
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_154
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_154 port map( A => S, Y => SB);
   UND1 : ND2_462 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_461 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_460 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_153 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_153;

architecture SYN_STRUCTURAL of MUX21_153 is

   component ND2_457
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_458
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_459
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_153
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_153 port map( A => S, Y => SB);
   UND1 : ND2_459 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_458 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_457 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_152 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_152;

architecture SYN_STRUCTURAL of MUX21_152 is

   component ND2_454
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_455
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_456
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_152
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_152 port map( A => S, Y => SB);
   UND1 : ND2_456 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_455 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_454 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_151 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_151;

architecture SYN_STRUCTURAL of MUX21_151 is

   component ND2_451
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_452
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_453
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_151
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_151 port map( A => S, Y => SB);
   UND1 : ND2_453 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_452 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_451 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_150 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_150;

architecture SYN_STRUCTURAL of MUX21_150 is

   component ND2_448
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_449
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_450
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_150
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_150 port map( A => S, Y => SB);
   UND1 : ND2_450 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_449 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_448 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_149 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_149;

architecture SYN_STRUCTURAL of MUX21_149 is

   component ND2_445
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_446
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_447
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_149
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_149 port map( A => S, Y => SB);
   UND1 : ND2_447 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_446 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_445 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_148 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_148;

architecture SYN_STRUCTURAL of MUX21_148 is

   component ND2_442
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_443
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_444
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_148
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_148 port map( A => S, Y => SB);
   UND1 : ND2_444 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_443 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_442 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_147 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_147;

architecture SYN_STRUCTURAL of MUX21_147 is

   component ND2_439
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_440
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_441
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_147
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_147 port map( A => S, Y => SB);
   UND1 : ND2_441 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_440 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_439 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_146 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_146;

architecture SYN_STRUCTURAL of MUX21_146 is

   component ND2_436
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_437
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_438
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_146
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_146 port map( A => S, Y => SB);
   UND1 : ND2_438 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_437 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_436 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_145 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_145;

architecture SYN_STRUCTURAL of MUX21_145 is

   component ND2_433
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_434
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_435
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_145
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_145 port map( A => S, Y => SB);
   UND1 : ND2_435 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_434 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_433 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_144 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_144;

architecture SYN_STRUCTURAL of MUX21_144 is

   component ND2_430
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_431
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_432
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_144
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_144 port map( A => S, Y => SB);
   UND1 : ND2_432 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_431 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_430 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_143 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_143;

architecture SYN_STRUCTURAL of MUX21_143 is

   component ND2_427
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_428
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_429
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_143
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_143 port map( A => S, Y => SB);
   UND1 : ND2_429 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_428 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_427 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_142 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_142;

architecture SYN_STRUCTURAL of MUX21_142 is

   component ND2_424
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_425
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_426
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_142
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_142 port map( A => S, Y => SB);
   UND1 : ND2_426 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_425 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_424 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_141 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_141;

architecture SYN_STRUCTURAL of MUX21_141 is

   component ND2_421
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_422
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_423
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_141
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_141 port map( A => S, Y => SB);
   UND1 : ND2_423 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_422 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_421 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_140 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_140;

architecture SYN_STRUCTURAL of MUX21_140 is

   component ND2_418
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_419
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_420
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_140
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_140 port map( A => S, Y => SB);
   UND1 : ND2_420 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_419 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_418 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_139 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_139;

architecture SYN_STRUCTURAL of MUX21_139 is

   component ND2_415
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_416
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_417
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_139
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_139 port map( A => S, Y => SB);
   UND1 : ND2_417 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_416 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_415 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_138 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_138;

architecture SYN_STRUCTURAL of MUX21_138 is

   component ND2_412
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_413
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_414
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_138
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_138 port map( A => S, Y => SB);
   UND1 : ND2_414 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_413 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_412 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_137 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_137;

architecture SYN_STRUCTURAL of MUX21_137 is

   component ND2_409
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_410
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_411
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_137
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_137 port map( A => S, Y => SB);
   UND1 : ND2_411 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_410 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_409 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_136 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_136;

architecture SYN_STRUCTURAL of MUX21_136 is

   component ND2_406
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_407
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_408
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_136
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_136 port map( A => S, Y => SB);
   UND1 : ND2_408 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_407 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_406 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_135 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_135;

architecture SYN_STRUCTURAL of MUX21_135 is

   component ND2_403
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_404
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_405
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_135
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_135 port map( A => S, Y => SB);
   UND1 : ND2_405 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_404 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_403 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_134 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_134;

architecture SYN_STRUCTURAL of MUX21_134 is

   component ND2_400
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_401
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_402
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_134
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_134 port map( A => S, Y => SB);
   UND1 : ND2_402 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_401 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_400 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_133 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_133;

architecture SYN_STRUCTURAL of MUX21_133 is

   component ND2_397
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_398
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_399
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_133
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_133 port map( A => S, Y => SB);
   UND1 : ND2_399 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_398 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_397 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_132 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_132;

architecture SYN_STRUCTURAL of MUX21_132 is

   component ND2_394
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_395
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_396
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_132
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_132 port map( A => S, Y => SB);
   UND1 : ND2_396 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_395 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_394 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_131 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_131;

architecture SYN_STRUCTURAL of MUX21_131 is

   component ND2_391
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_392
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_393
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_131
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_131 port map( A => S, Y => SB);
   UND1 : ND2_393 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_392 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_391 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_130 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_130;

architecture SYN_STRUCTURAL of MUX21_130 is

   component ND2_388
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_389
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_390
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_130
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_130 port map( A => S, Y => SB);
   UND1 : ND2_390 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_389 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_388 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_129 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_129;

architecture SYN_STRUCTURAL of MUX21_129 is

   component ND2_385
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_386
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_387
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_129
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_129 port map( A => S, Y => SB);
   UND1 : ND2_387 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_386 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_385 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_128 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_128;

architecture SYN_STRUCTURAL of MUX21_128 is

   component ND2_382
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_383
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_384
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_128
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_128 port map( A => S, Y => SB);
   UND1 : ND2_384 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_383 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_382 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_127 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_127;

architecture SYN_STRUCTURAL of MUX21_127 is

   component ND2_379
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_380
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_381
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_127
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_127 port map( A => S, Y => SB);
   UND1 : ND2_381 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_380 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_379 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_126 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_126;

architecture SYN_STRUCTURAL of MUX21_126 is

   component ND2_376
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_377
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_378
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_126
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_126 port map( A => S, Y => SB);
   UND1 : ND2_378 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_377 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_376 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_125 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_125;

architecture SYN_STRUCTURAL of MUX21_125 is

   component ND2_373
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_374
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_375
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_125
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_125 port map( A => S, Y => SB);
   UND1 : ND2_375 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_374 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_373 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_124 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_124;

architecture SYN_STRUCTURAL of MUX21_124 is

   component ND2_370
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_371
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_372
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_124
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_124 port map( A => S, Y => SB);
   UND1 : ND2_372 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_371 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_370 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_123 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_123;

architecture SYN_STRUCTURAL of MUX21_123 is

   component ND2_367
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_368
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_369
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_123
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_123 port map( A => S, Y => SB);
   UND1 : ND2_369 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_368 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_367 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_122 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_122;

architecture SYN_STRUCTURAL of MUX21_122 is

   component ND2_364
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_365
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_366
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_122
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_122 port map( A => S, Y => SB);
   UND1 : ND2_366 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_365 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_364 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_121 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_121;

architecture SYN_STRUCTURAL of MUX21_121 is

   component ND2_361
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_362
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_363
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_121
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_121 port map( A => S, Y => SB);
   UND1 : ND2_363 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_362 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_361 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_120 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_120;

architecture SYN_STRUCTURAL of MUX21_120 is

   component ND2_358
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_359
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_360
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_120
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_120 port map( A => S, Y => SB);
   UND1 : ND2_360 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_359 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_358 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_119 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_119;

architecture SYN_STRUCTURAL of MUX21_119 is

   component ND2_355
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_356
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_357
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_119
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_119 port map( A => S, Y => SB);
   UND1 : ND2_357 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_356 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_355 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_118 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_118;

architecture SYN_STRUCTURAL of MUX21_118 is

   component ND2_352
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_353
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_354
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_118
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_118 port map( A => S, Y => SB);
   UND1 : ND2_354 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_353 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_352 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_117 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_117;

architecture SYN_STRUCTURAL of MUX21_117 is

   component ND2_349
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_350
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_351
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_117
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_117 port map( A => S, Y => SB);
   UND1 : ND2_351 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_350 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_349 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_116 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_116;

architecture SYN_STRUCTURAL of MUX21_116 is

   component ND2_346
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_347
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_348
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_116
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_116 port map( A => S, Y => SB);
   UND1 : ND2_348 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_347 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_346 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_115 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_115;

architecture SYN_STRUCTURAL of MUX21_115 is

   component ND2_343
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_344
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_345
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_115
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_115 port map( A => S, Y => SB);
   UND1 : ND2_345 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_344 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_343 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_114 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_114;

architecture SYN_STRUCTURAL of MUX21_114 is

   component ND2_340
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_341
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_342
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_114
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_114 port map( A => S, Y => SB);
   UND1 : ND2_342 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_341 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_340 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_113 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_113;

architecture SYN_STRUCTURAL of MUX21_113 is

   component ND2_337
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_338
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_339
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_113
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_113 port map( A => S, Y => SB);
   UND1 : ND2_339 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_338 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_337 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_112 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_112;

architecture SYN_STRUCTURAL of MUX21_112 is

   component ND2_334
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_335
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_336
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_112
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_112 port map( A => S, Y => SB);
   UND1 : ND2_336 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_335 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_334 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_111 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_111;

architecture SYN_STRUCTURAL of MUX21_111 is

   component ND2_331
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_332
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_333
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_111
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_111 port map( A => S, Y => SB);
   UND1 : ND2_333 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_332 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_331 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_110 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_110;

architecture SYN_STRUCTURAL of MUX21_110 is

   component ND2_328
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_329
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_330
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_110
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_110 port map( A => S, Y => SB);
   UND1 : ND2_330 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_329 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_328 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_109 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_109;

architecture SYN_STRUCTURAL of MUX21_109 is

   component ND2_325
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_326
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_327
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_109
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_109 port map( A => S, Y => SB);
   UND1 : ND2_327 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_326 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_325 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_108 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_108;

architecture SYN_STRUCTURAL of MUX21_108 is

   component ND2_322
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_323
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_324
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_108
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_108 port map( A => S, Y => SB);
   UND1 : ND2_324 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_323 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_322 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_107 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_107;

architecture SYN_STRUCTURAL of MUX21_107 is

   component ND2_319
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_320
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_321
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_107
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_107 port map( A => S, Y => SB);
   UND1 : ND2_321 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_320 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_319 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_106 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_106;

architecture SYN_STRUCTURAL of MUX21_106 is

   component ND2_316
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_317
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_318
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_106
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_106 port map( A => S, Y => SB);
   UND1 : ND2_318 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_317 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_316 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_105 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_105;

architecture SYN_STRUCTURAL of MUX21_105 is

   component ND2_313
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_314
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_315
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_105
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_105 port map( A => S, Y => SB);
   UND1 : ND2_315 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_314 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_313 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_104 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_104;

architecture SYN_STRUCTURAL of MUX21_104 is

   component ND2_310
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_311
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_312
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_104
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_104 port map( A => S, Y => SB);
   UND1 : ND2_312 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_311 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_310 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_103 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_103;

architecture SYN_STRUCTURAL of MUX21_103 is

   component ND2_307
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_308
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_309
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_103
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_103 port map( A => S, Y => SB);
   UND1 : ND2_309 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_308 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_307 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_102 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_102;

architecture SYN_STRUCTURAL of MUX21_102 is

   component ND2_304
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_305
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_306
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_102
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_102 port map( A => S, Y => SB);
   UND1 : ND2_306 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_305 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_304 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_101 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_101;

architecture SYN_STRUCTURAL of MUX21_101 is

   component ND2_301
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_302
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_303
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_101
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_101 port map( A => S, Y => SB);
   UND1 : ND2_303 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_302 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_301 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_100 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_100;

architecture SYN_STRUCTURAL of MUX21_100 is

   component ND2_298
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_299
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_300
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_100
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_100 port map( A => S, Y => SB);
   UND1 : ND2_300 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_299 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_298 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_99 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_99;

architecture SYN_STRUCTURAL of MUX21_99 is

   component ND2_295
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_296
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_297
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_99
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_99 port map( A => S, Y => SB);
   UND1 : ND2_297 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_296 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_295 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_98 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_98;

architecture SYN_STRUCTURAL of MUX21_98 is

   component ND2_292
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_293
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_294
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_98
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_98 port map( A => S, Y => SB);
   UND1 : ND2_294 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_293 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_292 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_97 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_97;

architecture SYN_STRUCTURAL of MUX21_97 is

   component ND2_289
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_290
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_291
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_97
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_97 port map( A => S, Y => SB);
   UND1 : ND2_291 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_290 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_289 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_96 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_96;

architecture SYN_STRUCTURAL of MUX21_96 is

   component ND2_286
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_287
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_288
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_96
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_96 port map( A => S, Y => SB);
   UND1 : ND2_288 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_287 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_286 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_95 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_95;

architecture SYN_STRUCTURAL of MUX21_95 is

   component ND2_283
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_284
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_285
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_95
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_95 port map( A => S, Y => SB);
   UND1 : ND2_285 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_284 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_283 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_94 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_94;

architecture SYN_STRUCTURAL of MUX21_94 is

   component ND2_280
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_281
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_282
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_94
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_94 port map( A => S, Y => SB);
   UND1 : ND2_282 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_281 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_280 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_93 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_93;

architecture SYN_STRUCTURAL of MUX21_93 is

   component ND2_277
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_278
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_279
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_93
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_93 port map( A => S, Y => SB);
   UND1 : ND2_279 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_278 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_277 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_92 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_92;

architecture SYN_STRUCTURAL of MUX21_92 is

   component ND2_274
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_275
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_276
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_92
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_92 port map( A => S, Y => SB);
   UND1 : ND2_276 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_275 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_274 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_91 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_91;

architecture SYN_STRUCTURAL of MUX21_91 is

   component ND2_271
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_272
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_273
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_91
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_91 port map( A => S, Y => SB);
   UND1 : ND2_273 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_272 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_271 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_90 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_90;

architecture SYN_STRUCTURAL of MUX21_90 is

   component ND2_268
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_269
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_270
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_90
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_90 port map( A => S, Y => SB);
   UND1 : ND2_270 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_269 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_268 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_89 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_89;

architecture SYN_STRUCTURAL of MUX21_89 is

   component ND2_265
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_266
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_267
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_89
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_89 port map( A => S, Y => SB);
   UND1 : ND2_267 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_266 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_265 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_88 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_88;

architecture SYN_STRUCTURAL of MUX21_88 is

   component ND2_262
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_263
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_264
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_88
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_88 port map( A => S, Y => SB);
   UND1 : ND2_264 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_263 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_262 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_87 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_87;

architecture SYN_STRUCTURAL of MUX21_87 is

   component ND2_259
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_260
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_261
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_87
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_87 port map( A => S, Y => SB);
   UND1 : ND2_261 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_260 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_259 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_86 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_86;

architecture SYN_STRUCTURAL of MUX21_86 is

   component ND2_256
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_257
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_258
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_86
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_86 port map( A => S, Y => SB);
   UND1 : ND2_258 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_257 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_256 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_85 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_85;

architecture SYN_STRUCTURAL of MUX21_85 is

   component ND2_253
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_254
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_255
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_85
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_85 port map( A => S, Y => SB);
   UND1 : ND2_255 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_254 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_253 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_84 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_84;

architecture SYN_STRUCTURAL of MUX21_84 is

   component ND2_250
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_251
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_252
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_84
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_84 port map( A => S, Y => SB);
   UND1 : ND2_252 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_251 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_250 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_83 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_83;

architecture SYN_STRUCTURAL of MUX21_83 is

   component ND2_247
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_248
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_249
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_83
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_83 port map( A => S, Y => SB);
   UND1 : ND2_249 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_248 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_247 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_82 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_82;

architecture SYN_STRUCTURAL of MUX21_82 is

   component ND2_244
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_245
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_246
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_82
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_82 port map( A => S, Y => SB);
   UND1 : ND2_246 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_245 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_244 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_81 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_81;

architecture SYN_STRUCTURAL of MUX21_81 is

   component ND2_241
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_242
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_243
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_81
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_81 port map( A => S, Y => SB);
   UND1 : ND2_243 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_242 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_241 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_80 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_80;

architecture SYN_STRUCTURAL of MUX21_80 is

   component ND2_238
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_239
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_240
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_80
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_80 port map( A => S, Y => SB);
   UND1 : ND2_240 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_239 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_238 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_79 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_79;

architecture SYN_STRUCTURAL of MUX21_79 is

   component ND2_235
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_236
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_237
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_79
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_79 port map( A => S, Y => SB);
   UND1 : ND2_237 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_236 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_235 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_78 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_78;

architecture SYN_STRUCTURAL of MUX21_78 is

   component ND2_232
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_233
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_234
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_78
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_78 port map( A => S, Y => SB);
   UND1 : ND2_234 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_233 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_232 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_77 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_77;

architecture SYN_STRUCTURAL of MUX21_77 is

   component ND2_229
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_230
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_231
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_77
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_77 port map( A => S, Y => SB);
   UND1 : ND2_231 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_230 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_229 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_76 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_76;

architecture SYN_STRUCTURAL of MUX21_76 is

   component ND2_226
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_227
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_228
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_76
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_76 port map( A => S, Y => SB);
   UND1 : ND2_228 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_227 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_226 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_75 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_75;

architecture SYN_STRUCTURAL of MUX21_75 is

   component ND2_223
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_224
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_225
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_75
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_75 port map( A => S, Y => SB);
   UND1 : ND2_225 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_224 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_223 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_74 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_74;

architecture SYN_STRUCTURAL of MUX21_74 is

   component ND2_220
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_221
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_222
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_74
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_74 port map( A => S, Y => SB);
   UND1 : ND2_222 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_221 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_220 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_73 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_73;

architecture SYN_STRUCTURAL of MUX21_73 is

   component ND2_217
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_218
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_219
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_73
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_73 port map( A => S, Y => SB);
   UND1 : ND2_219 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_218 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_217 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_72 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_72;

architecture SYN_STRUCTURAL of MUX21_72 is

   component ND2_214
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_215
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_216
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_72
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_72 port map( A => S, Y => SB);
   UND1 : ND2_216 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_215 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_214 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_71 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_71;

architecture SYN_STRUCTURAL of MUX21_71 is

   component ND2_211
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_212
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_213
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_71
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_71 port map( A => S, Y => SB);
   UND1 : ND2_213 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_212 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_211 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_70 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_70;

architecture SYN_STRUCTURAL of MUX21_70 is

   component ND2_208
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_209
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_210
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_70
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_70 port map( A => S, Y => SB);
   UND1 : ND2_210 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_209 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_208 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_69 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_69;

architecture SYN_STRUCTURAL of MUX21_69 is

   component ND2_205
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_206
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_207
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_69
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_69 port map( A => S, Y => SB);
   UND1 : ND2_207 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_206 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_205 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_68 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_68;

architecture SYN_STRUCTURAL of MUX21_68 is

   component ND2_202
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_203
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_204
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_68
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_68 port map( A => S, Y => SB);
   UND1 : ND2_204 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_203 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_202 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_67 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_67;

architecture SYN_STRUCTURAL of MUX21_67 is

   component ND2_199
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_200
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_201
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_67
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_67 port map( A => S, Y => SB);
   UND1 : ND2_201 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_200 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_199 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_66 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_66;

architecture SYN_STRUCTURAL of MUX21_66 is

   component ND2_196
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_197
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_198
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_66
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_66 port map( A => S, Y => SB);
   UND1 : ND2_198 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_197 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_196 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_65 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_65;

architecture SYN_STRUCTURAL of MUX21_65 is

   component ND2_193
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_194
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_195
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_65
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_65 port map( A => S, Y => SB);
   UND1 : ND2_195 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_194 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_193 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_64 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_64;

architecture SYN_STRUCTURAL of MUX21_64 is

   component ND2_190
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_191
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_192
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_64
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_64 port map( A => S, Y => SB);
   UND1 : ND2_192 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_191 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_190 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_63 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_63;

architecture SYN_STRUCTURAL of MUX21_63 is

   component ND2_187
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_188
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_189
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_63
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_63 port map( A => S, Y => SB);
   UND1 : ND2_189 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_188 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_187 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_62 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_62;

architecture SYN_STRUCTURAL of MUX21_62 is

   component ND2_184
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_185
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_186
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_62
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_62 port map( A => S, Y => SB);
   UND1 : ND2_186 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_185 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_184 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_61 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_61;

architecture SYN_STRUCTURAL of MUX21_61 is

   component ND2_181
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_182
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_183
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_61
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_61 port map( A => S, Y => SB);
   UND1 : ND2_183 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_182 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_181 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_60 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_60;

architecture SYN_STRUCTURAL of MUX21_60 is

   component ND2_178
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_179
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_180
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_60
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_60 port map( A => S, Y => SB);
   UND1 : ND2_180 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_179 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_178 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_59 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_59;

architecture SYN_STRUCTURAL of MUX21_59 is

   component ND2_175
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_176
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_177
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_59
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_59 port map( A => S, Y => SB);
   UND1 : ND2_177 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_176 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_175 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_58 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_58;

architecture SYN_STRUCTURAL of MUX21_58 is

   component ND2_172
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_173
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_174
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_58
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_58 port map( A => S, Y => SB);
   UND1 : ND2_174 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_173 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_172 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_57 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_57;

architecture SYN_STRUCTURAL of MUX21_57 is

   component ND2_169
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_170
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_171
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_57
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_57 port map( A => S, Y => SB);
   UND1 : ND2_171 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_170 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_169 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_56 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_56;

architecture SYN_STRUCTURAL of MUX21_56 is

   component ND2_166
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_167
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_168
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_56
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_56 port map( A => S, Y => SB);
   UND1 : ND2_168 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_167 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_166 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_55 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_55;

architecture SYN_STRUCTURAL of MUX21_55 is

   component ND2_163
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_164
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_165
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_55
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_55 port map( A => S, Y => SB);
   UND1 : ND2_165 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_164 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_163 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_54 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_54;

architecture SYN_STRUCTURAL of MUX21_54 is

   component ND2_160
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_161
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_162
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_54
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_54 port map( A => S, Y => SB);
   UND1 : ND2_162 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_161 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_160 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_53 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_53;

architecture SYN_STRUCTURAL of MUX21_53 is

   component ND2_157
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_158
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_159
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_53
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_53 port map( A => S, Y => SB);
   UND1 : ND2_159 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_158 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_157 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_52 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_52;

architecture SYN_STRUCTURAL of MUX21_52 is

   component ND2_154
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_155
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_156
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_52
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_52 port map( A => S, Y => SB);
   UND1 : ND2_156 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_155 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_154 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_51 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_51;

architecture SYN_STRUCTURAL of MUX21_51 is

   component ND2_151
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_152
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_153
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_51
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_51 port map( A => S, Y => SB);
   UND1 : ND2_153 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_152 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_151 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_50 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_50;

architecture SYN_STRUCTURAL of MUX21_50 is

   component ND2_148
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_149
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_150
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_50
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_50 port map( A => S, Y => SB);
   UND1 : ND2_150 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_149 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_148 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_49 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_49;

architecture SYN_STRUCTURAL of MUX21_49 is

   component ND2_145
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_146
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_147
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_49
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_49 port map( A => S, Y => SB);
   UND1 : ND2_147 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_146 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_145 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_48 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_48;

architecture SYN_STRUCTURAL of MUX21_48 is

   component ND2_142
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_143
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_144
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_48
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_48 port map( A => S, Y => SB);
   UND1 : ND2_144 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_143 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_142 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_47 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_47;

architecture SYN_STRUCTURAL of MUX21_47 is

   component ND2_139
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_140
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_141
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_47
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_47 port map( A => S, Y => SB);
   UND1 : ND2_141 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_140 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_139 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_46 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_46;

architecture SYN_STRUCTURAL of MUX21_46 is

   component ND2_136
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_137
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_138
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_46
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_46 port map( A => S, Y => SB);
   UND1 : ND2_138 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_137 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_136 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_45 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_45;

architecture SYN_STRUCTURAL of MUX21_45 is

   component ND2_133
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_134
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_135
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_45
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_45 port map( A => S, Y => SB);
   UND1 : ND2_135 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_134 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_133 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_44 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_44;

architecture SYN_STRUCTURAL of MUX21_44 is

   component ND2_130
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_131
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_132
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_44
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_44 port map( A => S, Y => SB);
   UND1 : ND2_132 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_131 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_130 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_43 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_43;

architecture SYN_STRUCTURAL of MUX21_43 is

   component ND2_127
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_128
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_129
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_43
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_43 port map( A => S, Y => SB);
   UND1 : ND2_129 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_128 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_127 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_42 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_42;

architecture SYN_STRUCTURAL of MUX21_42 is

   component ND2_124
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_125
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_126
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_42
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_42 port map( A => S, Y => SB);
   UND1 : ND2_126 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_125 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_124 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_41 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_41;

architecture SYN_STRUCTURAL of MUX21_41 is

   component ND2_121
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_122
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_123
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_41
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_41 port map( A => S, Y => SB);
   UND1 : ND2_123 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_122 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_121 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_40 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_40;

architecture SYN_STRUCTURAL of MUX21_40 is

   component ND2_118
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_119
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_120
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_40
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_40 port map( A => S, Y => SB);
   UND1 : ND2_120 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_119 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_118 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_39 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_39;

architecture SYN_STRUCTURAL of MUX21_39 is

   component ND2_115
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_116
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_117
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_39
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_39 port map( A => S, Y => SB);
   UND1 : ND2_117 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_116 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_115 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_38 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_38;

architecture SYN_STRUCTURAL of MUX21_38 is

   component ND2_112
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_113
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_114
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_38
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_38 port map( A => S, Y => SB);
   UND1 : ND2_114 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_113 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_112 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_37 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_37;

architecture SYN_STRUCTURAL of MUX21_37 is

   component ND2_109
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_110
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_111
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_37
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_37 port map( A => S, Y => SB);
   UND1 : ND2_111 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_110 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_109 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_36 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_36;

architecture SYN_STRUCTURAL of MUX21_36 is

   component ND2_106
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_107
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_108
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_36
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_36 port map( A => S, Y => SB);
   UND1 : ND2_108 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_107 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_106 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_35 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_35;

architecture SYN_STRUCTURAL of MUX21_35 is

   component ND2_103
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_104
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_105
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_35
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_35 port map( A => S, Y => SB);
   UND1 : ND2_105 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_104 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_103 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_34 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_34;

architecture SYN_STRUCTURAL of MUX21_34 is

   component ND2_100
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_101
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_102
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_34
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_34 port map( A => S, Y => SB);
   UND1 : ND2_102 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_101 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_100 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_33 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_33;

architecture SYN_STRUCTURAL of MUX21_33 is

   component ND2_97
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_98
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_99
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_33
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_33 port map( A => S, Y => SB);
   UND1 : ND2_99 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_98 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_97 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_32 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_32;

architecture SYN_STRUCTURAL of MUX21_32 is

   component ND2_94
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_95
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_96
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_32
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_32 port map( A => S, Y => SB);
   UND1 : ND2_96 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_95 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_94 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_31 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_31;

architecture SYN_STRUCTURAL of MUX21_31 is

   component ND2_91
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_92
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_93
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_31
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_31 port map( A => S, Y => SB);
   UND1 : ND2_93 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_92 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_91 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_30 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_30;

architecture SYN_STRUCTURAL of MUX21_30 is

   component ND2_88
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_89
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_90
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_30
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_30 port map( A => S, Y => SB);
   UND1 : ND2_90 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_89 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_88 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_29 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_29;

architecture SYN_STRUCTURAL of MUX21_29 is

   component ND2_85
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_86
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_87
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_29
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_29 port map( A => S, Y => SB);
   UND1 : ND2_87 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_86 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_85 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_28 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_28;

architecture SYN_STRUCTURAL of MUX21_28 is

   component ND2_82
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_83
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_84
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_28
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_28 port map( A => S, Y => SB);
   UND1 : ND2_84 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_83 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_82 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_27 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_27;

architecture SYN_STRUCTURAL of MUX21_27 is

   component ND2_79
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_80
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_81
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_27
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_27 port map( A => S, Y => SB);
   UND1 : ND2_81 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_80 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_79 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_26 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_26;

architecture SYN_STRUCTURAL of MUX21_26 is

   component ND2_76
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_77
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_78
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_26
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_26 port map( A => S, Y => SB);
   UND1 : ND2_78 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_77 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_76 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_25 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_25;

architecture SYN_STRUCTURAL of MUX21_25 is

   component ND2_73
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_74
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_75
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_25
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_25 port map( A => S, Y => SB);
   UND1 : ND2_75 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_74 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_73 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_24 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_24;

architecture SYN_STRUCTURAL of MUX21_24 is

   component ND2_70
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_71
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_72
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_24
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_24 port map( A => S, Y => SB);
   UND1 : ND2_72 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_71 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_70 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_23 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_23;

architecture SYN_STRUCTURAL of MUX21_23 is

   component ND2_67
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_68
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_69
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_23
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_23 port map( A => S, Y => SB);
   UND1 : ND2_69 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_68 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_67 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_22 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_22;

architecture SYN_STRUCTURAL of MUX21_22 is

   component ND2_64
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_65
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_66
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_22
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_22 port map( A => S, Y => SB);
   UND1 : ND2_66 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_65 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_64 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_21 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_21;

architecture SYN_STRUCTURAL of MUX21_21 is

   component ND2_61
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_62
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_63
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_21
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_21 port map( A => S, Y => SB);
   UND1 : ND2_63 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_62 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_61 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_20 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_20;

architecture SYN_STRUCTURAL of MUX21_20 is

   component ND2_58
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_59
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_60
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_20
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_20 port map( A => S, Y => SB);
   UND1 : ND2_60 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_59 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_58 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_19 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_19;

architecture SYN_STRUCTURAL of MUX21_19 is

   component ND2_55
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_56
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_57
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_19
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_19 port map( A => S, Y => SB);
   UND1 : ND2_57 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_56 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_55 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_18 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_18;

architecture SYN_STRUCTURAL of MUX21_18 is

   component ND2_52
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_53
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_54
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_18
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_18 port map( A => S, Y => SB);
   UND1 : ND2_54 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_53 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_52 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_17 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_17;

architecture SYN_STRUCTURAL of MUX21_17 is

   component ND2_49
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_50
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_51
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_17
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_17 port map( A => S, Y => SB);
   UND1 : ND2_51 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_50 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_49 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_16 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_16;

architecture SYN_STRUCTURAL of MUX21_16 is

   component ND2_46
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_47
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_48
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_16
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_16 port map( A => S, Y => SB);
   UND1 : ND2_48 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_47 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_46 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_15 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_15;

architecture SYN_STRUCTURAL of MUX21_15 is

   component ND2_43
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_44
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_45
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_15
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_15 port map( A => S, Y => SB);
   UND1 : ND2_45 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_44 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_43 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_14 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_14;

architecture SYN_STRUCTURAL of MUX21_14 is

   component ND2_40
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_41
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_42
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_14
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_14 port map( A => S, Y => SB);
   UND1 : ND2_42 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_41 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_40 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_13 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_13;

architecture SYN_STRUCTURAL of MUX21_13 is

   component ND2_37
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_38
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_39
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_13
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_13 port map( A => S, Y => SB);
   UND1 : ND2_39 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_38 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_37 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_12 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_12;

architecture SYN_STRUCTURAL of MUX21_12 is

   component ND2_34
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_35
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_36
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_12
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_12 port map( A => S, Y => SB);
   UND1 : ND2_36 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_35 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_34 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_11 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_11;

architecture SYN_STRUCTURAL of MUX21_11 is

   component ND2_31
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_32
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_33
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_11
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_11 port map( A => S, Y => SB);
   UND1 : ND2_33 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_32 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_31 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_10 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_10;

architecture SYN_STRUCTURAL of MUX21_10 is

   component ND2_28
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_29
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_30
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_10
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_10 port map( A => S, Y => SB);
   UND1 : ND2_30 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_29 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_28 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_9 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_9;

architecture SYN_STRUCTURAL of MUX21_9 is

   component ND2_25
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_26
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_27
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_9
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_9 port map( A => S, Y => SB);
   UND1 : ND2_27 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_26 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_25 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_8 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_8;

architecture SYN_STRUCTURAL of MUX21_8 is

   component ND2_22
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_23
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_24
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_8
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_8 port map( A => S, Y => SB);
   UND1 : ND2_24 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_23 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_22 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_7 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_7;

architecture SYN_STRUCTURAL of MUX21_7 is

   component ND2_19
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_20
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_21
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_7
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_7 port map( A => S, Y => SB);
   UND1 : ND2_21 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_20 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_19 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_6 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_6;

architecture SYN_STRUCTURAL of MUX21_6 is

   component ND2_16
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_17
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_18
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_6
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_6 port map( A => S, Y => SB);
   UND1 : ND2_18 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_17 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_16 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_5 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_5;

architecture SYN_STRUCTURAL of MUX21_5 is

   component ND2_13
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_14
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_15
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_5
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_5 port map( A => S, Y => SB);
   UND1 : ND2_15 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_14 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_13 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_4 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_4;

architecture SYN_STRUCTURAL of MUX21_4 is

   component ND2_10
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_11
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_12
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_4 port map( A => S, Y => SB);
   UND1 : ND2_12 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_11 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_10 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_3 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_3;

architecture SYN_STRUCTURAL of MUX21_3 is

   component ND2_7
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_8
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_9
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_3
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_3 port map( A => S, Y => SB);
   UND1 : ND2_9 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_8 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_7 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_2 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_2;

architecture SYN_STRUCTURAL of MUX21_2 is

   component ND2_4
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_5
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_6
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_2 port map( A => S, Y => SB);
   UND1 : ND2_6 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_5 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_4 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_1 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_1;

architecture SYN_STRUCTURAL of MUX21_1 is

   component ND2_1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_3
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_1 port map( A => S, Y => SB);
   UND1 : ND2_3 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_2 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_1 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity FA_47 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_47;

architecture SYN_Behavioural of FA_47 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => c_in, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => c_out);
   U3 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n1, B2 => c_in, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n1);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity FA_46 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_46;

architecture SYN_Behavioural of FA_46 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => c_in, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => c_out);
   U3 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n1, B2 => c_in, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n1);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity FA_45 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_45;

architecture SYN_Behavioural of FA_45 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => c_in, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => c_out);
   U3 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n1, B2 => c_in, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n1);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity FA_44 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_44;

architecture SYN_Behavioural of FA_44 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => c_in, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => c_out);
   U3 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n1, B2 => c_in, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n1);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity FA_43 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_43;

architecture SYN_Behavioural of FA_43 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => c_in, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => c_out);
   U3 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n1, B2 => c_in, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n1);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity FA_42 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_42;

architecture SYN_Behavioural of FA_42 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => c_in, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => c_out);
   U3 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n1, B2 => c_in, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n1);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity FA_41 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_41;

architecture SYN_Behavioural of FA_41 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => c_in, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => c_out);
   U3 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n1, B2 => c_in, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n1);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity FA_40 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_40;

architecture SYN_Behavioural of FA_40 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => c_in, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => c_out);
   U3 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n1, B2 => c_in, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n1);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity FA_39 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_39;

architecture SYN_Behavioural of FA_39 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => c_in, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => c_out);
   U3 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n1, B2 => c_in, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n1);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity FA_38 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_38;

architecture SYN_Behavioural of FA_38 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => c_in, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => c_out);
   U3 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n1, B2 => c_in, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n1);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity FA_37 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_37;

architecture SYN_Behavioural of FA_37 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => c_in, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => c_out);
   U3 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n1, B2 => c_in, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n1);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity FA_36 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_36;

architecture SYN_Behavioural of FA_36 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => c_in, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => c_out);
   U3 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n1, B2 => c_in, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n1);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity FA_35 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_35;

architecture SYN_Behavioural of FA_35 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => c_in, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => c_out);
   U3 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n1, B2 => c_in, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n1);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity FA_34 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_34;

architecture SYN_Behavioural of FA_34 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => c_in, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => c_out);
   U3 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n1, B2 => c_in, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n1);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity FA_33 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_33;

architecture SYN_Behavioural of FA_33 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => c_in, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => c_out);
   U3 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n1, B2 => c_in, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n1);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity FA_32 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_32;

architecture SYN_Behavioural of FA_32 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => c_in, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => c_out);
   U3 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n1, B2 => c_in, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n1);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity FA_31 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_31;

architecture SYN_Behavioural of FA_31 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => c_in, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => c_out);
   U3 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n1, B2 => c_in, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n1);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity FA_30 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_30;

architecture SYN_Behavioural of FA_30 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => c_in, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => c_out);
   U3 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n1, B2 => c_in, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n1);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity FA_29 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_29;

architecture SYN_Behavioural of FA_29 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => c_in, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => c_out);
   U3 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n1, B2 => c_in, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n1);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity FA_28 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_28;

architecture SYN_Behavioural of FA_28 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => c_in, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => c_out);
   U3 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n1, B2 => c_in, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n1);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity FA_27 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_27;

architecture SYN_Behavioural of FA_27 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => c_in, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => c_out);
   U3 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n1, B2 => c_in, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n1);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity FA_26 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_26;

architecture SYN_Behavioural of FA_26 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => c_in, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => c_out);
   U3 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n1, B2 => c_in, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n1);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity FA_25 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_25;

architecture SYN_Behavioural of FA_25 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => c_in, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => c_out);
   U3 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n1, B2 => c_in, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n1);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity FA_24 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_24;

architecture SYN_Behavioural of FA_24 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => c_in, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => c_out);
   U3 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n1, B2 => c_in, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n1);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity FA_23 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_23;

architecture SYN_Behavioural of FA_23 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => c_in, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => c_out);
   U3 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n1, B2 => c_in, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n1);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity FA_22 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_22;

architecture SYN_Behavioural of FA_22 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => c_in, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => c_out);
   U3 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n1, B2 => c_in, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n1);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity FA_21 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_21;

architecture SYN_Behavioural of FA_21 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => c_in, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => c_out);
   U3 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n1, B2 => c_in, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n1);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity FA_20 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_20;

architecture SYN_Behavioural of FA_20 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => c_in, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => c_out);
   U3 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n1, B2 => c_in, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n1);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity FA_19 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_19;

architecture SYN_Behavioural of FA_19 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => c_in, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => c_out);
   U3 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n1, B2 => c_in, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n1);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity FA_18 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_18;

architecture SYN_Behavioural of FA_18 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => c_in, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => c_out);
   U3 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n1, B2 => c_in, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n1);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity FA_17 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_17;

architecture SYN_Behavioural of FA_17 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => c_in, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => c_out);
   U3 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n1, B2 => c_in, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n1);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity FA_16 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_16;

architecture SYN_Behavioural of FA_16 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => c_in, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => c_out);
   U3 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n1, B2 => c_in, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n1);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity FA_15 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_15;

architecture SYN_Behavioural of FA_15 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => c_in, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => c_out);
   U3 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n1, B2 => c_in, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n1);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity FA_14 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_14;

architecture SYN_Behavioural of FA_14 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => c_in, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => c_out);
   U3 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n1, B2 => c_in, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n1);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity FA_13 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_13;

architecture SYN_Behavioural of FA_13 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => c_in, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => c_out);
   U3 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n1, B2 => c_in, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n1);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity FA_12 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_12;

architecture SYN_Behavioural of FA_12 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => c_in, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => c_out);
   U3 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n1, B2 => c_in, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n1);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity FA_11 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_11;

architecture SYN_Behavioural of FA_11 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => c_in, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => c_out);
   U3 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n1, B2 => c_in, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n1);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity FA_10 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_10;

architecture SYN_Behavioural of FA_10 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => c_in, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => c_out);
   U3 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n1, B2 => c_in, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n1);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity FA_9 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_9;

architecture SYN_Behavioural of FA_9 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => c_in, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => c_out);
   U3 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n1, B2 => c_in, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n1);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity FA_8 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_8;

architecture SYN_Behavioural of FA_8 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => c_in, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => c_out);
   U3 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n1, B2 => c_in, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n1);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity FA_7 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_7;

architecture SYN_Behavioural of FA_7 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => c_in, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => c_out);
   U3 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n1, B2 => c_in, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n1);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity FA_6 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_6;

architecture SYN_Behavioural of FA_6 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => c_in, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => c_out);
   U3 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n1, B2 => c_in, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n1);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity FA_5 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_5;

architecture SYN_Behavioural of FA_5 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => c_in, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => c_out);
   U3 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n1, B2 => c_in, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n1);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity FA_4 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_4;

architecture SYN_Behavioural of FA_4 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => c_in, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => c_out);
   U3 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n1, B2 => c_in, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n1);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity FA_3 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_3;

architecture SYN_Behavioural of FA_3 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => c_in, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => c_out);
   U3 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n1, B2 => c_in, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n1);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity FA_2 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_2;

architecture SYN_Behavioural of FA_2 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => c_in, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => c_out);
   U3 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n1, B2 => c_in, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n1);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity FA_1 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_1;

architecture SYN_Behavioural of FA_1 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => c_in, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => c_out);
   U3 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n1, B2 => c_in, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n1);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_GENERIC_NBIT16_15 is

   port( A, B : in std_logic_vector (15 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (15 downto 0));

end MUX21_GENERIC_NBIT16_15;

architecture SYN_STRUCTURAL of MUX21_GENERIC_NBIT16_15 is

   component MUX21_225
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_226
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_227
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_228
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_229
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_230
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_231
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_232
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_233
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_234
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_235
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_236
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_237
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_238
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_239
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_240
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUX21GENI_0 : MUX21_240 port map( A => A(0), B => B(0), S => SEL, Y => Y(0))
                           ;
   MUX21GENI_1 : MUX21_239 port map( A => A(1), B => B(1), S => SEL, Y => Y(1))
                           ;
   MUX21GENI_2 : MUX21_238 port map( A => A(2), B => B(2), S => SEL, Y => Y(2))
                           ;
   MUX21GENI_3 : MUX21_237 port map( A => A(3), B => B(3), S => SEL, Y => Y(3))
                           ;
   MUX21GENI_4 : MUX21_236 port map( A => A(4), B => B(4), S => SEL, Y => Y(4))
                           ;
   MUX21GENI_5 : MUX21_235 port map( A => A(5), B => B(5), S => SEL, Y => Y(5))
                           ;
   MUX21GENI_6 : MUX21_234 port map( A => A(6), B => B(6), S => SEL, Y => Y(6))
                           ;
   MUX21GENI_7 : MUX21_233 port map( A => A(7), B => B(7), S => SEL, Y => Y(7))
                           ;
   MUX21GENI_8 : MUX21_232 port map( A => A(8), B => B(8), S => SEL, Y => Y(8))
                           ;
   MUX21GENI_9 : MUX21_231 port map( A => A(9), B => B(9), S => SEL, Y => Y(9))
                           ;
   MUX21GENI_10 : MUX21_230 port map( A => A(10), B => B(10), S => SEL, Y => 
                           Y(10));
   MUX21GENI_11 : MUX21_229 port map( A => A(11), B => B(11), S => SEL, Y => 
                           Y(11));
   MUX21GENI_12 : MUX21_228 port map( A => A(12), B => B(12), S => SEL, Y => 
                           Y(12));
   MUX21GENI_13 : MUX21_227 port map( A => A(13), B => B(13), S => SEL, Y => 
                           Y(13));
   MUX21GENI_14 : MUX21_226 port map( A => A(14), B => B(14), S => SEL, Y => 
                           Y(14));
   MUX21GENI_15 : MUX21_225 port map( A => A(15), B => B(15), S => SEL, Y => 
                           Y(15));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_GENERIC_NBIT16_14 is

   port( A, B : in std_logic_vector (15 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (15 downto 0));

end MUX21_GENERIC_NBIT16_14;

architecture SYN_STRUCTURAL of MUX21_GENERIC_NBIT16_14 is

   component MUX21_209
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_210
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_211
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_212
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_213
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_214
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_215
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_216
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_217
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_218
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_219
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_220
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_221
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_222
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_223
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_224
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUX21GENI_0 : MUX21_224 port map( A => A(0), B => B(0), S => SEL, Y => Y(0))
                           ;
   MUX21GENI_1 : MUX21_223 port map( A => A(1), B => B(1), S => SEL, Y => Y(1))
                           ;
   MUX21GENI_2 : MUX21_222 port map( A => A(2), B => B(2), S => SEL, Y => Y(2))
                           ;
   MUX21GENI_3 : MUX21_221 port map( A => A(3), B => B(3), S => SEL, Y => Y(3))
                           ;
   MUX21GENI_4 : MUX21_220 port map( A => A(4), B => B(4), S => SEL, Y => Y(4))
                           ;
   MUX21GENI_5 : MUX21_219 port map( A => A(5), B => B(5), S => SEL, Y => Y(5))
                           ;
   MUX21GENI_6 : MUX21_218 port map( A => A(6), B => B(6), S => SEL, Y => Y(6))
                           ;
   MUX21GENI_7 : MUX21_217 port map( A => A(7), B => B(7), S => SEL, Y => Y(7))
                           ;
   MUX21GENI_8 : MUX21_216 port map( A => A(8), B => B(8), S => SEL, Y => Y(8))
                           ;
   MUX21GENI_9 : MUX21_215 port map( A => A(9), B => B(9), S => SEL, Y => Y(9))
                           ;
   MUX21GENI_10 : MUX21_214 port map( A => A(10), B => B(10), S => SEL, Y => 
                           Y(10));
   MUX21GENI_11 : MUX21_213 port map( A => A(11), B => B(11), S => SEL, Y => 
                           Y(11));
   MUX21GENI_12 : MUX21_212 port map( A => A(12), B => B(12), S => SEL, Y => 
                           Y(12));
   MUX21GENI_13 : MUX21_211 port map( A => A(13), B => B(13), S => SEL, Y => 
                           Y(13));
   MUX21GENI_14 : MUX21_210 port map( A => A(14), B => B(14), S => SEL, Y => 
                           Y(14));
   MUX21GENI_15 : MUX21_209 port map( A => A(15), B => B(15), S => SEL, Y => 
                           Y(15));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_GENERIC_NBIT16_13 is

   port( A, B : in std_logic_vector (15 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (15 downto 0));

end MUX21_GENERIC_NBIT16_13;

architecture SYN_STRUCTURAL of MUX21_GENERIC_NBIT16_13 is

   component MUX21_193
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_194
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_195
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_196
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_197
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_198
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_199
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_200
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_201
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_202
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_203
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_204
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_205
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_206
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_207
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_208
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUX21GENI_0 : MUX21_208 port map( A => A(0), B => B(0), S => SEL, Y => Y(0))
                           ;
   MUX21GENI_1 : MUX21_207 port map( A => A(1), B => B(1), S => SEL, Y => Y(1))
                           ;
   MUX21GENI_2 : MUX21_206 port map( A => A(2), B => B(2), S => SEL, Y => Y(2))
                           ;
   MUX21GENI_3 : MUX21_205 port map( A => A(3), B => B(3), S => SEL, Y => Y(3))
                           ;
   MUX21GENI_4 : MUX21_204 port map( A => A(4), B => B(4), S => SEL, Y => Y(4))
                           ;
   MUX21GENI_5 : MUX21_203 port map( A => A(5), B => B(5), S => SEL, Y => Y(5))
                           ;
   MUX21GENI_6 : MUX21_202 port map( A => A(6), B => B(6), S => SEL, Y => Y(6))
                           ;
   MUX21GENI_7 : MUX21_201 port map( A => A(7), B => B(7), S => SEL, Y => Y(7))
                           ;
   MUX21GENI_8 : MUX21_200 port map( A => A(8), B => B(8), S => SEL, Y => Y(8))
                           ;
   MUX21GENI_9 : MUX21_199 port map( A => A(9), B => B(9), S => SEL, Y => Y(9))
                           ;
   MUX21GENI_10 : MUX21_198 port map( A => A(10), B => B(10), S => SEL, Y => 
                           Y(10));
   MUX21GENI_11 : MUX21_197 port map( A => A(11), B => B(11), S => SEL, Y => 
                           Y(11));
   MUX21GENI_12 : MUX21_196 port map( A => A(12), B => B(12), S => SEL, Y => 
                           Y(12));
   MUX21GENI_13 : MUX21_195 port map( A => A(13), B => B(13), S => SEL, Y => 
                           Y(13));
   MUX21GENI_14 : MUX21_194 port map( A => A(14), B => B(14), S => SEL, Y => 
                           Y(14));
   MUX21GENI_15 : MUX21_193 port map( A => A(15), B => B(15), S => SEL, Y => 
                           Y(15));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_GENERIC_NBIT16_12 is

   port( A, B : in std_logic_vector (15 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (15 downto 0));

end MUX21_GENERIC_NBIT16_12;

architecture SYN_STRUCTURAL of MUX21_GENERIC_NBIT16_12 is

   component MUX21_177
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_178
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_179
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_180
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_181
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_182
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_183
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_184
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_185
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_186
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_187
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_188
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_189
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_190
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_191
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_192
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUX21GENI_0 : MUX21_192 port map( A => A(0), B => B(0), S => SEL, Y => Y(0))
                           ;
   MUX21GENI_1 : MUX21_191 port map( A => A(1), B => B(1), S => SEL, Y => Y(1))
                           ;
   MUX21GENI_2 : MUX21_190 port map( A => A(2), B => B(2), S => SEL, Y => Y(2))
                           ;
   MUX21GENI_3 : MUX21_189 port map( A => A(3), B => B(3), S => SEL, Y => Y(3))
                           ;
   MUX21GENI_4 : MUX21_188 port map( A => A(4), B => B(4), S => SEL, Y => Y(4))
                           ;
   MUX21GENI_5 : MUX21_187 port map( A => A(5), B => B(5), S => SEL, Y => Y(5))
                           ;
   MUX21GENI_6 : MUX21_186 port map( A => A(6), B => B(6), S => SEL, Y => Y(6))
                           ;
   MUX21GENI_7 : MUX21_185 port map( A => A(7), B => B(7), S => SEL, Y => Y(7))
                           ;
   MUX21GENI_8 : MUX21_184 port map( A => A(8), B => B(8), S => SEL, Y => Y(8))
                           ;
   MUX21GENI_9 : MUX21_183 port map( A => A(9), B => B(9), S => SEL, Y => Y(9))
                           ;
   MUX21GENI_10 : MUX21_182 port map( A => A(10), B => B(10), S => SEL, Y => 
                           Y(10));
   MUX21GENI_11 : MUX21_181 port map( A => A(11), B => B(11), S => SEL, Y => 
                           Y(11));
   MUX21GENI_12 : MUX21_180 port map( A => A(12), B => B(12), S => SEL, Y => 
                           Y(12));
   MUX21GENI_13 : MUX21_179 port map( A => A(13), B => B(13), S => SEL, Y => 
                           Y(13));
   MUX21GENI_14 : MUX21_178 port map( A => A(14), B => B(14), S => SEL, Y => 
                           Y(14));
   MUX21GENI_15 : MUX21_177 port map( A => A(15), B => B(15), S => SEL, Y => 
                           Y(15));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_GENERIC_NBIT16_11 is

   port( A, B : in std_logic_vector (15 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (15 downto 0));

end MUX21_GENERIC_NBIT16_11;

architecture SYN_STRUCTURAL of MUX21_GENERIC_NBIT16_11 is

   component MUX21_161
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_162
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_163
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_164
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_165
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_166
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_167
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_168
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_169
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_170
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_171
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_172
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_173
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_174
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_175
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_176
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUX21GENI_0 : MUX21_176 port map( A => A(0), B => B(0), S => SEL, Y => Y(0))
                           ;
   MUX21GENI_1 : MUX21_175 port map( A => A(1), B => B(1), S => SEL, Y => Y(1))
                           ;
   MUX21GENI_2 : MUX21_174 port map( A => A(2), B => B(2), S => SEL, Y => Y(2))
                           ;
   MUX21GENI_3 : MUX21_173 port map( A => A(3), B => B(3), S => SEL, Y => Y(3))
                           ;
   MUX21GENI_4 : MUX21_172 port map( A => A(4), B => B(4), S => SEL, Y => Y(4))
                           ;
   MUX21GENI_5 : MUX21_171 port map( A => A(5), B => B(5), S => SEL, Y => Y(5))
                           ;
   MUX21GENI_6 : MUX21_170 port map( A => A(6), B => B(6), S => SEL, Y => Y(6))
                           ;
   MUX21GENI_7 : MUX21_169 port map( A => A(7), B => B(7), S => SEL, Y => Y(7))
                           ;
   MUX21GENI_8 : MUX21_168 port map( A => A(8), B => B(8), S => SEL, Y => Y(8))
                           ;
   MUX21GENI_9 : MUX21_167 port map( A => A(9), B => B(9), S => SEL, Y => Y(9))
                           ;
   MUX21GENI_10 : MUX21_166 port map( A => A(10), B => B(10), S => SEL, Y => 
                           Y(10));
   MUX21GENI_11 : MUX21_165 port map( A => A(11), B => B(11), S => SEL, Y => 
                           Y(11));
   MUX21GENI_12 : MUX21_164 port map( A => A(12), B => B(12), S => SEL, Y => 
                           Y(12));
   MUX21GENI_13 : MUX21_163 port map( A => A(13), B => B(13), S => SEL, Y => 
                           Y(13));
   MUX21GENI_14 : MUX21_162 port map( A => A(14), B => B(14), S => SEL, Y => 
                           Y(14));
   MUX21GENI_15 : MUX21_161 port map( A => A(15), B => B(15), S => SEL, Y => 
                           Y(15));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_GENERIC_NBIT16_10 is

   port( A, B : in std_logic_vector (15 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (15 downto 0));

end MUX21_GENERIC_NBIT16_10;

architecture SYN_STRUCTURAL of MUX21_GENERIC_NBIT16_10 is

   component MUX21_145
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_146
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_147
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_148
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_149
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_150
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_151
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_152
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_153
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_154
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_155
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_156
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_157
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_158
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_159
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_160
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUX21GENI_0 : MUX21_160 port map( A => A(0), B => B(0), S => SEL, Y => Y(0))
                           ;
   MUX21GENI_1 : MUX21_159 port map( A => A(1), B => B(1), S => SEL, Y => Y(1))
                           ;
   MUX21GENI_2 : MUX21_158 port map( A => A(2), B => B(2), S => SEL, Y => Y(2))
                           ;
   MUX21GENI_3 : MUX21_157 port map( A => A(3), B => B(3), S => SEL, Y => Y(3))
                           ;
   MUX21GENI_4 : MUX21_156 port map( A => A(4), B => B(4), S => SEL, Y => Y(4))
                           ;
   MUX21GENI_5 : MUX21_155 port map( A => A(5), B => B(5), S => SEL, Y => Y(5))
                           ;
   MUX21GENI_6 : MUX21_154 port map( A => A(6), B => B(6), S => SEL, Y => Y(6))
                           ;
   MUX21GENI_7 : MUX21_153 port map( A => A(7), B => B(7), S => SEL, Y => Y(7))
                           ;
   MUX21GENI_8 : MUX21_152 port map( A => A(8), B => B(8), S => SEL, Y => Y(8))
                           ;
   MUX21GENI_9 : MUX21_151 port map( A => A(9), B => B(9), S => SEL, Y => Y(9))
                           ;
   MUX21GENI_10 : MUX21_150 port map( A => A(10), B => B(10), S => SEL, Y => 
                           Y(10));
   MUX21GENI_11 : MUX21_149 port map( A => A(11), B => B(11), S => SEL, Y => 
                           Y(11));
   MUX21GENI_12 : MUX21_148 port map( A => A(12), B => B(12), S => SEL, Y => 
                           Y(12));
   MUX21GENI_13 : MUX21_147 port map( A => A(13), B => B(13), S => SEL, Y => 
                           Y(13));
   MUX21GENI_14 : MUX21_146 port map( A => A(14), B => B(14), S => SEL, Y => 
                           Y(14));
   MUX21GENI_15 : MUX21_145 port map( A => A(15), B => B(15), S => SEL, Y => 
                           Y(15));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_GENERIC_NBIT16_9 is

   port( A, B : in std_logic_vector (15 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (15 downto 0));

end MUX21_GENERIC_NBIT16_9;

architecture SYN_STRUCTURAL of MUX21_GENERIC_NBIT16_9 is

   component MUX21_129
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_130
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_131
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_132
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_133
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_134
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_135
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_136
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_137
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_138
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_139
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_140
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_141
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_142
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_143
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_144
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUX21GENI_0 : MUX21_144 port map( A => A(0), B => B(0), S => SEL, Y => Y(0))
                           ;
   MUX21GENI_1 : MUX21_143 port map( A => A(1), B => B(1), S => SEL, Y => Y(1))
                           ;
   MUX21GENI_2 : MUX21_142 port map( A => A(2), B => B(2), S => SEL, Y => Y(2))
                           ;
   MUX21GENI_3 : MUX21_141 port map( A => A(3), B => B(3), S => SEL, Y => Y(3))
                           ;
   MUX21GENI_4 : MUX21_140 port map( A => A(4), B => B(4), S => SEL, Y => Y(4))
                           ;
   MUX21GENI_5 : MUX21_139 port map( A => A(5), B => B(5), S => SEL, Y => Y(5))
                           ;
   MUX21GENI_6 : MUX21_138 port map( A => A(6), B => B(6), S => SEL, Y => Y(6))
                           ;
   MUX21GENI_7 : MUX21_137 port map( A => A(7), B => B(7), S => SEL, Y => Y(7))
                           ;
   MUX21GENI_8 : MUX21_136 port map( A => A(8), B => B(8), S => SEL, Y => Y(8))
                           ;
   MUX21GENI_9 : MUX21_135 port map( A => A(9), B => B(9), S => SEL, Y => Y(9))
                           ;
   MUX21GENI_10 : MUX21_134 port map( A => A(10), B => B(10), S => SEL, Y => 
                           Y(10));
   MUX21GENI_11 : MUX21_133 port map( A => A(11), B => B(11), S => SEL, Y => 
                           Y(11));
   MUX21GENI_12 : MUX21_132 port map( A => A(12), B => B(12), S => SEL, Y => 
                           Y(12));
   MUX21GENI_13 : MUX21_131 port map( A => A(13), B => B(13), S => SEL, Y => 
                           Y(13));
   MUX21GENI_14 : MUX21_130 port map( A => A(14), B => B(14), S => SEL, Y => 
                           Y(14));
   MUX21GENI_15 : MUX21_129 port map( A => A(15), B => B(15), S => SEL, Y => 
                           Y(15));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_GENERIC_NBIT16_8 is

   port( A, B : in std_logic_vector (15 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (15 downto 0));

end MUX21_GENERIC_NBIT16_8;

architecture SYN_STRUCTURAL of MUX21_GENERIC_NBIT16_8 is

   component MUX21_113
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_114
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_115
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_116
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_117
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_118
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_119
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_120
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_121
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_122
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_123
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_124
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_125
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_126
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_127
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_128
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUX21GENI_0 : MUX21_128 port map( A => A(0), B => B(0), S => SEL, Y => Y(0))
                           ;
   MUX21GENI_1 : MUX21_127 port map( A => A(1), B => B(1), S => SEL, Y => Y(1))
                           ;
   MUX21GENI_2 : MUX21_126 port map( A => A(2), B => B(2), S => SEL, Y => Y(2))
                           ;
   MUX21GENI_3 : MUX21_125 port map( A => A(3), B => B(3), S => SEL, Y => Y(3))
                           ;
   MUX21GENI_4 : MUX21_124 port map( A => A(4), B => B(4), S => SEL, Y => Y(4))
                           ;
   MUX21GENI_5 : MUX21_123 port map( A => A(5), B => B(5), S => SEL, Y => Y(5))
                           ;
   MUX21GENI_6 : MUX21_122 port map( A => A(6), B => B(6), S => SEL, Y => Y(6))
                           ;
   MUX21GENI_7 : MUX21_121 port map( A => A(7), B => B(7), S => SEL, Y => Y(7))
                           ;
   MUX21GENI_8 : MUX21_120 port map( A => A(8), B => B(8), S => SEL, Y => Y(8))
                           ;
   MUX21GENI_9 : MUX21_119 port map( A => A(9), B => B(9), S => SEL, Y => Y(9))
                           ;
   MUX21GENI_10 : MUX21_118 port map( A => A(10), B => B(10), S => SEL, Y => 
                           Y(10));
   MUX21GENI_11 : MUX21_117 port map( A => A(11), B => B(11), S => SEL, Y => 
                           Y(11));
   MUX21GENI_12 : MUX21_116 port map( A => A(12), B => B(12), S => SEL, Y => 
                           Y(12));
   MUX21GENI_13 : MUX21_115 port map( A => A(13), B => B(13), S => SEL, Y => 
                           Y(13));
   MUX21GENI_14 : MUX21_114 port map( A => A(14), B => B(14), S => SEL, Y => 
                           Y(14));
   MUX21GENI_15 : MUX21_113 port map( A => A(15), B => B(15), S => SEL, Y => 
                           Y(15));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_GENERIC_NBIT16_7 is

   port( A, B : in std_logic_vector (15 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (15 downto 0));

end MUX21_GENERIC_NBIT16_7;

architecture SYN_STRUCTURAL of MUX21_GENERIC_NBIT16_7 is

   component MUX21_97
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_98
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_99
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_100
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_101
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_102
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_103
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_104
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_105
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_106
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_107
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_108
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_109
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_110
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_111
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_112
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUX21GENI_0 : MUX21_112 port map( A => A(0), B => B(0), S => SEL, Y => Y(0))
                           ;
   MUX21GENI_1 : MUX21_111 port map( A => A(1), B => B(1), S => SEL, Y => Y(1))
                           ;
   MUX21GENI_2 : MUX21_110 port map( A => A(2), B => B(2), S => SEL, Y => Y(2))
                           ;
   MUX21GENI_3 : MUX21_109 port map( A => A(3), B => B(3), S => SEL, Y => Y(3))
                           ;
   MUX21GENI_4 : MUX21_108 port map( A => A(4), B => B(4), S => SEL, Y => Y(4))
                           ;
   MUX21GENI_5 : MUX21_107 port map( A => A(5), B => B(5), S => SEL, Y => Y(5))
                           ;
   MUX21GENI_6 : MUX21_106 port map( A => A(6), B => B(6), S => SEL, Y => Y(6))
                           ;
   MUX21GENI_7 : MUX21_105 port map( A => A(7), B => B(7), S => SEL, Y => Y(7))
                           ;
   MUX21GENI_8 : MUX21_104 port map( A => A(8), B => B(8), S => SEL, Y => Y(8))
                           ;
   MUX21GENI_9 : MUX21_103 port map( A => A(9), B => B(9), S => SEL, Y => Y(9))
                           ;
   MUX21GENI_10 : MUX21_102 port map( A => A(10), B => B(10), S => SEL, Y => 
                           Y(10));
   MUX21GENI_11 : MUX21_101 port map( A => A(11), B => B(11), S => SEL, Y => 
                           Y(11));
   MUX21GENI_12 : MUX21_100 port map( A => A(12), B => B(12), S => SEL, Y => 
                           Y(12));
   MUX21GENI_13 : MUX21_99 port map( A => A(13), B => B(13), S => SEL, Y => 
                           Y(13));
   MUX21GENI_14 : MUX21_98 port map( A => A(14), B => B(14), S => SEL, Y => 
                           Y(14));
   MUX21GENI_15 : MUX21_97 port map( A => A(15), B => B(15), S => SEL, Y => 
                           Y(15));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_GENERIC_NBIT16_6 is

   port( A, B : in std_logic_vector (15 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (15 downto 0));

end MUX21_GENERIC_NBIT16_6;

architecture SYN_STRUCTURAL of MUX21_GENERIC_NBIT16_6 is

   component MUX21_81
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_82
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_83
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_84
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_85
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_86
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_87
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_88
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_89
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_90
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_91
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_92
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_93
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_94
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_95
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_96
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUX21GENI_0 : MUX21_96 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUX21GENI_1 : MUX21_95 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUX21GENI_2 : MUX21_94 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUX21GENI_3 : MUX21_93 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));
   MUX21GENI_4 : MUX21_92 port map( A => A(4), B => B(4), S => SEL, Y => Y(4));
   MUX21GENI_5 : MUX21_91 port map( A => A(5), B => B(5), S => SEL, Y => Y(5));
   MUX21GENI_6 : MUX21_90 port map( A => A(6), B => B(6), S => SEL, Y => Y(6));
   MUX21GENI_7 : MUX21_89 port map( A => A(7), B => B(7), S => SEL, Y => Y(7));
   MUX21GENI_8 : MUX21_88 port map( A => A(8), B => B(8), S => SEL, Y => Y(8));
   MUX21GENI_9 : MUX21_87 port map( A => A(9), B => B(9), S => SEL, Y => Y(9));
   MUX21GENI_10 : MUX21_86 port map( A => A(10), B => B(10), S => SEL, Y => 
                           Y(10));
   MUX21GENI_11 : MUX21_85 port map( A => A(11), B => B(11), S => SEL, Y => 
                           Y(11));
   MUX21GENI_12 : MUX21_84 port map( A => A(12), B => B(12), S => SEL, Y => 
                           Y(12));
   MUX21GENI_13 : MUX21_83 port map( A => A(13), B => B(13), S => SEL, Y => 
                           Y(13));
   MUX21GENI_14 : MUX21_82 port map( A => A(14), B => B(14), S => SEL, Y => 
                           Y(14));
   MUX21GENI_15 : MUX21_81 port map( A => A(15), B => B(15), S => SEL, Y => 
                           Y(15));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_GENERIC_NBIT16_5 is

   port( A, B : in std_logic_vector (15 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (15 downto 0));

end MUX21_GENERIC_NBIT16_5;

architecture SYN_STRUCTURAL of MUX21_GENERIC_NBIT16_5 is

   component MUX21_65
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_66
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_67
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_68
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_69
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_70
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_71
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_72
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_73
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_74
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_75
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_76
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_77
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_78
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_79
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_80
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUX21GENI_0 : MUX21_80 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUX21GENI_1 : MUX21_79 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUX21GENI_2 : MUX21_78 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUX21GENI_3 : MUX21_77 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));
   MUX21GENI_4 : MUX21_76 port map( A => A(4), B => B(4), S => SEL, Y => Y(4));
   MUX21GENI_5 : MUX21_75 port map( A => A(5), B => B(5), S => SEL, Y => Y(5));
   MUX21GENI_6 : MUX21_74 port map( A => A(6), B => B(6), S => SEL, Y => Y(6));
   MUX21GENI_7 : MUX21_73 port map( A => A(7), B => B(7), S => SEL, Y => Y(7));
   MUX21GENI_8 : MUX21_72 port map( A => A(8), B => B(8), S => SEL, Y => Y(8));
   MUX21GENI_9 : MUX21_71 port map( A => A(9), B => B(9), S => SEL, Y => Y(9));
   MUX21GENI_10 : MUX21_70 port map( A => A(10), B => B(10), S => SEL, Y => 
                           Y(10));
   MUX21GENI_11 : MUX21_69 port map( A => A(11), B => B(11), S => SEL, Y => 
                           Y(11));
   MUX21GENI_12 : MUX21_68 port map( A => A(12), B => B(12), S => SEL, Y => 
                           Y(12));
   MUX21GENI_13 : MUX21_67 port map( A => A(13), B => B(13), S => SEL, Y => 
                           Y(13));
   MUX21GENI_14 : MUX21_66 port map( A => A(14), B => B(14), S => SEL, Y => 
                           Y(14));
   MUX21GENI_15 : MUX21_65 port map( A => A(15), B => B(15), S => SEL, Y => 
                           Y(15));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_GENERIC_NBIT16_4 is

   port( A, B : in std_logic_vector (15 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (15 downto 0));

end MUX21_GENERIC_NBIT16_4;

architecture SYN_STRUCTURAL of MUX21_GENERIC_NBIT16_4 is

   component MUX21_49
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_50
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_51
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_52
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_53
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_54
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_55
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_56
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_57
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_58
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_59
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_60
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_61
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_62
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_63
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_64
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUX21GENI_0 : MUX21_64 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUX21GENI_1 : MUX21_63 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUX21GENI_2 : MUX21_62 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUX21GENI_3 : MUX21_61 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));
   MUX21GENI_4 : MUX21_60 port map( A => A(4), B => B(4), S => SEL, Y => Y(4));
   MUX21GENI_5 : MUX21_59 port map( A => A(5), B => B(5), S => SEL, Y => Y(5));
   MUX21GENI_6 : MUX21_58 port map( A => A(6), B => B(6), S => SEL, Y => Y(6));
   MUX21GENI_7 : MUX21_57 port map( A => A(7), B => B(7), S => SEL, Y => Y(7));
   MUX21GENI_8 : MUX21_56 port map( A => A(8), B => B(8), S => SEL, Y => Y(8));
   MUX21GENI_9 : MUX21_55 port map( A => A(9), B => B(9), S => SEL, Y => Y(9));
   MUX21GENI_10 : MUX21_54 port map( A => A(10), B => B(10), S => SEL, Y => 
                           Y(10));
   MUX21GENI_11 : MUX21_53 port map( A => A(11), B => B(11), S => SEL, Y => 
                           Y(11));
   MUX21GENI_12 : MUX21_52 port map( A => A(12), B => B(12), S => SEL, Y => 
                           Y(12));
   MUX21GENI_13 : MUX21_51 port map( A => A(13), B => B(13), S => SEL, Y => 
                           Y(13));
   MUX21GENI_14 : MUX21_50 port map( A => A(14), B => B(14), S => SEL, Y => 
                           Y(14));
   MUX21GENI_15 : MUX21_49 port map( A => A(15), B => B(15), S => SEL, Y => 
                           Y(15));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_GENERIC_NBIT16_3 is

   port( A, B : in std_logic_vector (15 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (15 downto 0));

end MUX21_GENERIC_NBIT16_3;

architecture SYN_STRUCTURAL of MUX21_GENERIC_NBIT16_3 is

   component MUX21_33
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_34
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_35
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_36
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_37
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_38
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_39
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_40
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_41
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_42
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_43
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_44
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_45
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_46
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_47
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_48
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUX21GENI_0 : MUX21_48 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUX21GENI_1 : MUX21_47 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUX21GENI_2 : MUX21_46 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUX21GENI_3 : MUX21_45 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));
   MUX21GENI_4 : MUX21_44 port map( A => A(4), B => B(4), S => SEL, Y => Y(4));
   MUX21GENI_5 : MUX21_43 port map( A => A(5), B => B(5), S => SEL, Y => Y(5));
   MUX21GENI_6 : MUX21_42 port map( A => A(6), B => B(6), S => SEL, Y => Y(6));
   MUX21GENI_7 : MUX21_41 port map( A => A(7), B => B(7), S => SEL, Y => Y(7));
   MUX21GENI_8 : MUX21_40 port map( A => A(8), B => B(8), S => SEL, Y => Y(8));
   MUX21GENI_9 : MUX21_39 port map( A => A(9), B => B(9), S => SEL, Y => Y(9));
   MUX21GENI_10 : MUX21_38 port map( A => A(10), B => B(10), S => SEL, Y => 
                           Y(10));
   MUX21GENI_11 : MUX21_37 port map( A => A(11), B => B(11), S => SEL, Y => 
                           Y(11));
   MUX21GENI_12 : MUX21_36 port map( A => A(12), B => B(12), S => SEL, Y => 
                           Y(12));
   MUX21GENI_13 : MUX21_35 port map( A => A(13), B => B(13), S => SEL, Y => 
                           Y(13));
   MUX21GENI_14 : MUX21_34 port map( A => A(14), B => B(14), S => SEL, Y => 
                           Y(14));
   MUX21GENI_15 : MUX21_33 port map( A => A(15), B => B(15), S => SEL, Y => 
                           Y(15));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_GENERIC_NBIT16_2 is

   port( A, B : in std_logic_vector (15 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (15 downto 0));

end MUX21_GENERIC_NBIT16_2;

architecture SYN_STRUCTURAL of MUX21_GENERIC_NBIT16_2 is

   component MUX21_17
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_18
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_19
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_20
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_21
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_22
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_23
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_24
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_25
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_26
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_27
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_28
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_29
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_30
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_31
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_32
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUX21GENI_0 : MUX21_32 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUX21GENI_1 : MUX21_31 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUX21GENI_2 : MUX21_30 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUX21GENI_3 : MUX21_29 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));
   MUX21GENI_4 : MUX21_28 port map( A => A(4), B => B(4), S => SEL, Y => Y(4));
   MUX21GENI_5 : MUX21_27 port map( A => A(5), B => B(5), S => SEL, Y => Y(5));
   MUX21GENI_6 : MUX21_26 port map( A => A(6), B => B(6), S => SEL, Y => Y(6));
   MUX21GENI_7 : MUX21_25 port map( A => A(7), B => B(7), S => SEL, Y => Y(7));
   MUX21GENI_8 : MUX21_24 port map( A => A(8), B => B(8), S => SEL, Y => Y(8));
   MUX21GENI_9 : MUX21_23 port map( A => A(9), B => B(9), S => SEL, Y => Y(9));
   MUX21GENI_10 : MUX21_22 port map( A => A(10), B => B(10), S => SEL, Y => 
                           Y(10));
   MUX21GENI_11 : MUX21_21 port map( A => A(11), B => B(11), S => SEL, Y => 
                           Y(11));
   MUX21GENI_12 : MUX21_20 port map( A => A(12), B => B(12), S => SEL, Y => 
                           Y(12));
   MUX21GENI_13 : MUX21_19 port map( A => A(13), B => B(13), S => SEL, Y => 
                           Y(13));
   MUX21GENI_14 : MUX21_18 port map( A => A(14), B => B(14), S => SEL, Y => 
                           Y(14));
   MUX21GENI_15 : MUX21_17 port map( A => A(15), B => B(15), S => SEL, Y => 
                           Y(15));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_GENERIC_NBIT16_1 is

   port( A, B : in std_logic_vector (15 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (15 downto 0));

end MUX21_GENERIC_NBIT16_1;

architecture SYN_STRUCTURAL of MUX21_GENERIC_NBIT16_1 is

   component MUX21_1
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_2
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_3
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_4
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_5
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_6
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_7
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_8
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_9
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_10
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_11
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_12
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_13
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_14
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_15
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_16
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUX21GENI_0 : MUX21_16 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUX21GENI_1 : MUX21_15 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUX21GENI_2 : MUX21_14 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUX21GENI_3 : MUX21_13 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));
   MUX21GENI_4 : MUX21_12 port map( A => A(4), B => B(4), S => SEL, Y => Y(4));
   MUX21GENI_5 : MUX21_11 port map( A => A(5), B => B(5), S => SEL, Y => Y(5));
   MUX21GENI_6 : MUX21_10 port map( A => A(6), B => B(6), S => SEL, Y => Y(6));
   MUX21GENI_7 : MUX21_9 port map( A => A(7), B => B(7), S => SEL, Y => Y(7));
   MUX21GENI_8 : MUX21_8 port map( A => A(8), B => B(8), S => SEL, Y => Y(8));
   MUX21GENI_9 : MUX21_7 port map( A => A(9), B => B(9), S => SEL, Y => Y(9));
   MUX21GENI_10 : MUX21_6 port map( A => A(10), B => B(10), S => SEL, Y => 
                           Y(10));
   MUX21GENI_11 : MUX21_5 port map( A => A(11), B => B(11), S => SEL, Y => 
                           Y(11));
   MUX21GENI_12 : MUX21_4 port map( A => A(12), B => B(12), S => SEL, Y => 
                           Y(12));
   MUX21GENI_13 : MUX21_3 port map( A => A(13), B => B(13), S => SEL, Y => 
                           Y(13));
   MUX21GENI_14 : MUX21_2 port map( A => A(14), B => B(14), S => SEL, Y => 
                           Y(14));
   MUX21GENI_15 : MUX21_1 port map( A => A(15), B => B(15), S => SEL, Y => 
                           Y(15));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity RCA_size16_2 is

   port( a, b : in std_logic_vector (15 downto 0);  c_in : in std_logic;  c_out
         : out std_logic;  sum : out std_logic_vector (15 downto 0));

end RCA_size16_2;

architecture SYN_Structural of RCA_size16_2 is

   component FA_17
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_18
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_19
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_20
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_21
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_22
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_23
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_24
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_25
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_26
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_27
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_28
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_29
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_30
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_31
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_32
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   signal temp_15_port, temp_14_port, temp_13_port, temp_12_port, temp_11_port,
      temp_10_port, temp_9_port, temp_8_port, temp_7_port, temp_6_port, 
      temp_5_port, temp_4_port, temp_3_port, temp_2_port, temp_1_port : 
      std_logic;

begin
   
   fa_i_0 : FA_32 port map( a => a(0), b => b(0), c_in => c_in, c_out => 
                           temp_1_port, s => sum(0));
   fa_i_1 : FA_31 port map( a => a(1), b => b(1), c_in => temp_1_port, c_out =>
                           temp_2_port, s => sum(1));
   fa_i_2 : FA_30 port map( a => a(2), b => b(2), c_in => temp_2_port, c_out =>
                           temp_3_port, s => sum(2));
   fa_i_3 : FA_29 port map( a => a(3), b => b(3), c_in => temp_3_port, c_out =>
                           temp_4_port, s => sum(3));
   fa_i_4 : FA_28 port map( a => a(4), b => b(4), c_in => temp_4_port, c_out =>
                           temp_5_port, s => sum(4));
   fa_i_5 : FA_27 port map( a => a(5), b => b(5), c_in => temp_5_port, c_out =>
                           temp_6_port, s => sum(5));
   fa_i_6 : FA_26 port map( a => a(6), b => b(6), c_in => temp_6_port, c_out =>
                           temp_7_port, s => sum(6));
   fa_i_7 : FA_25 port map( a => a(7), b => b(7), c_in => temp_7_port, c_out =>
                           temp_8_port, s => sum(7));
   fa_i_8 : FA_24 port map( a => a(8), b => b(8), c_in => temp_8_port, c_out =>
                           temp_9_port, s => sum(8));
   fa_i_9 : FA_23 port map( a => a(9), b => b(9), c_in => temp_9_port, c_out =>
                           temp_10_port, s => sum(9));
   fa_i_10 : FA_22 port map( a => a(10), b => b(10), c_in => temp_10_port, 
                           c_out => temp_11_port, s => sum(10));
   fa_i_11 : FA_21 port map( a => a(11), b => b(11), c_in => temp_11_port, 
                           c_out => temp_12_port, s => sum(11));
   fa_i_12 : FA_20 port map( a => a(12), b => b(12), c_in => temp_12_port, 
                           c_out => temp_13_port, s => sum(12));
   fa_i_13 : FA_19 port map( a => a(13), b => b(13), c_in => temp_13_port, 
                           c_out => temp_14_port, s => sum(13));
   fa_i_14 : FA_18 port map( a => a(14), b => b(14), c_in => temp_14_port, 
                           c_out => temp_15_port, s => sum(14));
   fa_i_15 : FA_17 port map( a => a(15), b => b(15), c_in => temp_15_port, 
                           c_out => c_out, s => sum(15));

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity RCA_size16_1 is

   port( a, b : in std_logic_vector (15 downto 0);  c_in : in std_logic;  c_out
         : out std_logic;  sum : out std_logic_vector (15 downto 0));

end RCA_size16_1;

architecture SYN_Structural of RCA_size16_1 is

   component FA_1
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_2
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_3
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_4
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_5
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_6
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_7
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_8
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_9
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_10
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_11
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_12
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_13
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_14
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_15
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_16
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   signal temp_15_port, temp_14_port, temp_13_port, temp_12_port, temp_11_port,
      temp_10_port, temp_9_port, temp_8_port, temp_7_port, temp_6_port, 
      temp_5_port, temp_4_port, temp_3_port, temp_2_port, temp_1_port : 
      std_logic;

begin
   
   fa_i_0 : FA_16 port map( a => a(0), b => b(0), c_in => c_in, c_out => 
                           temp_1_port, s => sum(0));
   fa_i_1 : FA_15 port map( a => a(1), b => b(1), c_in => temp_1_port, c_out =>
                           temp_2_port, s => sum(1));
   fa_i_2 : FA_14 port map( a => a(2), b => b(2), c_in => temp_2_port, c_out =>
                           temp_3_port, s => sum(2));
   fa_i_3 : FA_13 port map( a => a(3), b => b(3), c_in => temp_3_port, c_out =>
                           temp_4_port, s => sum(3));
   fa_i_4 : FA_12 port map( a => a(4), b => b(4), c_in => temp_4_port, c_out =>
                           temp_5_port, s => sum(4));
   fa_i_5 : FA_11 port map( a => a(5), b => b(5), c_in => temp_5_port, c_out =>
                           temp_6_port, s => sum(5));
   fa_i_6 : FA_10 port map( a => a(6), b => b(6), c_in => temp_6_port, c_out =>
                           temp_7_port, s => sum(6));
   fa_i_7 : FA_9 port map( a => a(7), b => b(7), c_in => temp_7_port, c_out => 
                           temp_8_port, s => sum(7));
   fa_i_8 : FA_8 port map( a => a(8), b => b(8), c_in => temp_8_port, c_out => 
                           temp_9_port, s => sum(8));
   fa_i_9 : FA_7 port map( a => a(9), b => b(9), c_in => temp_9_port, c_out => 
                           temp_10_port, s => sum(9));
   fa_i_10 : FA_6 port map( a => a(10), b => b(10), c_in => temp_10_port, c_out
                           => temp_11_port, s => sum(10));
   fa_i_11 : FA_5 port map( a => a(11), b => b(11), c_in => temp_11_port, c_out
                           => temp_12_port, s => sum(11));
   fa_i_12 : FA_4 port map( a => a(12), b => b(12), c_in => temp_12_port, c_out
                           => temp_13_port, s => sum(12));
   fa_i_13 : FA_3 port map( a => a(13), b => b(13), c_in => temp_13_port, c_out
                           => temp_14_port, s => sum(13));
   fa_i_14 : FA_2 port map( a => a(14), b => b(14), c_in => temp_14_port, c_out
                           => temp_15_port, s => sum(14));
   fa_i_15 : FA_1 port map( a => a(15), b => b(15), c_in => temp_15_port, c_out
                           => c_out, s => sum(15));

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX51_GENERIC_NBIT16_3 is

   port( A0, A1, A2, A3, A4 : in std_logic_vector (15 downto 0);  SEL : in 
         std_logic_vector (2 downto 0);  Y : out std_logic_vector (15 downto 0)
         );

end MUX51_GENERIC_NBIT16_3;

architecture SYN_STRUCTURAL of MUX51_GENERIC_NBIT16_3 is

   component MUX21_GENERIC_NBIT16_9
      port( A, B : in std_logic_vector (15 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (15 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT16_10
      port( A, B : in std_logic_vector (15 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (15 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT16_11
      port( A, B : in std_logic_vector (15 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (15 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT16_12
      port( A, B : in std_logic_vector (15 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (15 downto 0));
   end component;
   
   signal Y0_15_port, Y0_14_port, Y0_13_port, Y0_12_port, Y0_11_port, 
      Y0_10_port, Y0_9_port, Y0_8_port, Y0_7_port, Y0_6_port, Y0_5_port, 
      Y0_4_port, Y0_3_port, Y0_2_port, Y0_1_port, Y0_0_port, Y1_15_port, 
      Y1_14_port, Y1_13_port, Y1_12_port, Y1_11_port, Y1_10_port, Y1_9_port, 
      Y1_8_port, Y1_7_port, Y1_6_port, Y1_5_port, Y1_4_port, Y1_3_port, 
      Y1_2_port, Y1_1_port, Y1_0_port, Y2_15_port, Y2_14_port, Y2_13_port, 
      Y2_12_port, Y2_11_port, Y2_10_port, Y2_9_port, Y2_8_port, Y2_7_port, 
      Y2_6_port, Y2_5_port, Y2_4_port, Y2_3_port, Y2_2_port, Y2_1_port, 
      Y2_0_port : std_logic;

begin
   
   mux000 : MUX21_GENERIC_NBIT16_12 port map( A(15) => A0(15), A(14) => A0(14),
                           A(13) => A0(13), A(12) => A0(12), A(11) => A0(11), 
                           A(10) => A0(10), A(9) => A0(9), A(8) => A0(8), A(7) 
                           => A0(7), A(6) => A0(6), A(5) => A0(5), A(4) => 
                           A0(4), A(3) => A0(3), A(2) => A0(2), A(1) => A0(1), 
                           A(0) => A0(0), B(15) => A1(15), B(14) => A1(14), 
                           B(13) => A1(13), B(12) => A1(12), B(11) => A1(11), 
                           B(10) => A1(10), B(9) => A1(9), B(8) => A1(8), B(7) 
                           => A1(7), B(6) => A1(6), B(5) => A1(5), B(4) => 
                           A1(4), B(3) => A1(3), B(2) => A1(2), B(1) => A1(1), 
                           B(0) => A1(0), SEL => SEL(2), Y(15) => Y0_15_port, 
                           Y(14) => Y0_14_port, Y(13) => Y0_13_port, Y(12) => 
                           Y0_12_port, Y(11) => Y0_11_port, Y(10) => Y0_10_port
                           , Y(9) => Y0_9_port, Y(8) => Y0_8_port, Y(7) => 
                           Y0_7_port, Y(6) => Y0_6_port, Y(5) => Y0_5_port, 
                           Y(4) => Y0_4_port, Y(3) => Y0_3_port, Y(2) => 
                           Y0_2_port, Y(1) => Y0_1_port, Y(0) => Y0_0_port);
   mux100 : MUX21_GENERIC_NBIT16_11 port map( A(15) => A2(15), A(14) => A2(14),
                           A(13) => A2(13), A(12) => A2(12), A(11) => A2(11), 
                           A(10) => A2(10), A(9) => A2(9), A(8) => A2(8), A(7) 
                           => A2(7), A(6) => A2(6), A(5) => A2(5), A(4) => 
                           A2(4), A(3) => A2(3), A(2) => A2(2), A(1) => A2(1), 
                           A(0) => A2(0), B(15) => A3(15), B(14) => A3(14), 
                           B(13) => A3(13), B(12) => A3(12), B(11) => A3(11), 
                           B(10) => A3(10), B(9) => A3(9), B(8) => A3(8), B(7) 
                           => A3(7), B(6) => A3(6), B(5) => A3(5), B(4) => 
                           A3(4), B(3) => A3(3), B(2) => A3(2), B(1) => A3(1), 
                           B(0) => A3(0), SEL => SEL(2), Y(15) => Y1_15_port, 
                           Y(14) => Y1_14_port, Y(13) => Y1_13_port, Y(12) => 
                           Y1_12_port, Y(11) => Y1_11_port, Y(10) => Y1_10_port
                           , Y(9) => Y1_9_port, Y(8) => Y1_8_port, Y(7) => 
                           Y1_7_port, Y(6) => Y1_6_port, Y(5) => Y1_5_port, 
                           Y(4) => Y1_4_port, Y(3) => Y1_3_port, Y(2) => 
                           Y1_2_port, Y(1) => Y1_1_port, Y(0) => Y1_0_port);
   mux010 : MUX21_GENERIC_NBIT16_10 port map( A(15) => Y0_15_port, A(14) => 
                           Y0_14_port, A(13) => Y0_13_port, A(12) => Y0_12_port
                           , A(11) => Y0_11_port, A(10) => Y0_10_port, A(9) => 
                           Y0_9_port, A(8) => Y0_8_port, A(7) => Y0_7_port, 
                           A(6) => Y0_6_port, A(5) => Y0_5_port, A(4) => 
                           Y0_4_port, A(3) => Y0_3_port, A(2) => Y0_2_port, 
                           A(1) => Y0_1_port, A(0) => Y0_0_port, B(15) => 
                           Y1_15_port, B(14) => Y1_14_port, B(13) => Y1_13_port
                           , B(12) => Y1_12_port, B(11) => Y1_11_port, B(10) =>
                           Y1_10_port, B(9) => Y1_9_port, B(8) => Y1_8_port, 
                           B(7) => Y1_7_port, B(6) => Y1_6_port, B(5) => 
                           Y1_5_port, B(4) => Y1_4_port, B(3) => Y1_3_port, 
                           B(2) => Y1_2_port, B(1) => Y1_1_port, B(0) => 
                           Y1_0_port, SEL => SEL(1), Y(15) => Y2_15_port, Y(14)
                           => Y2_14_port, Y(13) => Y2_13_port, Y(12) => 
                           Y2_12_port, Y(11) => Y2_11_port, Y(10) => Y2_10_port
                           , Y(9) => Y2_9_port, Y(8) => Y2_8_port, Y(7) => 
                           Y2_7_port, Y(6) => Y2_6_port, Y(5) => Y2_5_port, 
                           Y(4) => Y2_4_port, Y(3) => Y2_3_port, Y(2) => 
                           Y2_2_port, Y(1) => Y2_1_port, Y(0) => Y2_0_port);
   mux001 : MUX21_GENERIC_NBIT16_9 port map( A(15) => Y2_15_port, A(14) => 
                           Y2_14_port, A(13) => Y2_13_port, A(12) => Y2_12_port
                           , A(11) => Y2_11_port, A(10) => Y2_10_port, A(9) => 
                           Y2_9_port, A(8) => Y2_8_port, A(7) => Y2_7_port, 
                           A(6) => Y2_6_port, A(5) => Y2_5_port, A(4) => 
                           Y2_4_port, A(3) => Y2_3_port, A(2) => Y2_2_port, 
                           A(1) => Y2_1_port, A(0) => Y2_0_port, B(15) => 
                           A4(15), B(14) => A4(14), B(13) => A4(13), B(12) => 
                           A4(12), B(11) => A4(11), B(10) => A4(10), B(9) => 
                           A4(9), B(8) => A4(8), B(7) => A4(7), B(6) => A4(6), 
                           B(5) => A4(5), B(4) => A4(4), B(3) => A4(3), B(2) =>
                           A4(2), B(1) => A4(1), B(0) => A4(0), SEL => SEL(0), 
                           Y(15) => Y(15), Y(14) => Y(14), Y(13) => Y(13), 
                           Y(12) => Y(12), Y(11) => Y(11), Y(10) => Y(10), Y(9)
                           => Y(9), Y(8) => Y(8), Y(7) => Y(7), Y(6) => Y(6), 
                           Y(5) => Y(5), Y(4) => Y(4), Y(3) => Y(3), Y(2) => 
                           Y(2), Y(1) => Y(1), Y(0) => Y(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX51_GENERIC_NBIT16_2 is

   port( A0, A1, A2, A3, A4 : in std_logic_vector (15 downto 0);  SEL : in 
         std_logic_vector (2 downto 0);  Y : out std_logic_vector (15 downto 0)
         );

end MUX51_GENERIC_NBIT16_2;

architecture SYN_STRUCTURAL of MUX51_GENERIC_NBIT16_2 is

   component MUX21_GENERIC_NBIT16_5
      port( A, B : in std_logic_vector (15 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (15 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT16_6
      port( A, B : in std_logic_vector (15 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (15 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT16_7
      port( A, B : in std_logic_vector (15 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (15 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT16_8
      port( A, B : in std_logic_vector (15 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (15 downto 0));
   end component;
   
   signal Y0_15_port, Y0_14_port, Y0_13_port, Y0_12_port, Y0_11_port, 
      Y0_10_port, Y0_9_port, Y0_8_port, Y0_7_port, Y0_6_port, Y0_5_port, 
      Y0_4_port, Y0_3_port, Y0_2_port, Y0_1_port, Y0_0_port, Y1_15_port, 
      Y1_14_port, Y1_13_port, Y1_12_port, Y1_11_port, Y1_10_port, Y1_9_port, 
      Y1_8_port, Y1_7_port, Y1_6_port, Y1_5_port, Y1_4_port, Y1_3_port, 
      Y1_2_port, Y1_1_port, Y1_0_port, Y2_15_port, Y2_14_port, Y2_13_port, 
      Y2_12_port, Y2_11_port, Y2_10_port, Y2_9_port, Y2_8_port, Y2_7_port, 
      Y2_6_port, Y2_5_port, Y2_4_port, Y2_3_port, Y2_2_port, Y2_1_port, 
      Y2_0_port : std_logic;

begin
   
   mux000 : MUX21_GENERIC_NBIT16_8 port map( A(15) => A0(15), A(14) => A0(14), 
                           A(13) => A0(13), A(12) => A0(12), A(11) => A0(11), 
                           A(10) => A0(10), A(9) => A0(9), A(8) => A0(8), A(7) 
                           => A0(7), A(6) => A0(6), A(5) => A0(5), A(4) => 
                           A0(4), A(3) => A0(3), A(2) => A0(2), A(1) => A0(1), 
                           A(0) => A0(0), B(15) => A1(15), B(14) => A1(14), 
                           B(13) => A1(13), B(12) => A1(12), B(11) => A1(11), 
                           B(10) => A1(10), B(9) => A1(9), B(8) => A1(8), B(7) 
                           => A1(7), B(6) => A1(6), B(5) => A1(5), B(4) => 
                           A1(4), B(3) => A1(3), B(2) => A1(2), B(1) => A1(1), 
                           B(0) => A1(0), SEL => SEL(2), Y(15) => Y0_15_port, 
                           Y(14) => Y0_14_port, Y(13) => Y0_13_port, Y(12) => 
                           Y0_12_port, Y(11) => Y0_11_port, Y(10) => Y0_10_port
                           , Y(9) => Y0_9_port, Y(8) => Y0_8_port, Y(7) => 
                           Y0_7_port, Y(6) => Y0_6_port, Y(5) => Y0_5_port, 
                           Y(4) => Y0_4_port, Y(3) => Y0_3_port, Y(2) => 
                           Y0_2_port, Y(1) => Y0_1_port, Y(0) => Y0_0_port);
   mux100 : MUX21_GENERIC_NBIT16_7 port map( A(15) => A2(15), A(14) => A2(14), 
                           A(13) => A2(13), A(12) => A2(12), A(11) => A2(11), 
                           A(10) => A2(10), A(9) => A2(9), A(8) => A2(8), A(7) 
                           => A2(7), A(6) => A2(6), A(5) => A2(5), A(4) => 
                           A2(4), A(3) => A2(3), A(2) => A2(2), A(1) => A2(1), 
                           A(0) => A2(0), B(15) => A3(15), B(14) => A3(14), 
                           B(13) => A3(13), B(12) => A3(12), B(11) => A3(11), 
                           B(10) => A3(10), B(9) => A3(9), B(8) => A3(8), B(7) 
                           => A3(7), B(6) => A3(6), B(5) => A3(5), B(4) => 
                           A3(4), B(3) => A3(3), B(2) => A3(2), B(1) => A3(1), 
                           B(0) => A3(0), SEL => SEL(2), Y(15) => Y1_15_port, 
                           Y(14) => Y1_14_port, Y(13) => Y1_13_port, Y(12) => 
                           Y1_12_port, Y(11) => Y1_11_port, Y(10) => Y1_10_port
                           , Y(9) => Y1_9_port, Y(8) => Y1_8_port, Y(7) => 
                           Y1_7_port, Y(6) => Y1_6_port, Y(5) => Y1_5_port, 
                           Y(4) => Y1_4_port, Y(3) => Y1_3_port, Y(2) => 
                           Y1_2_port, Y(1) => Y1_1_port, Y(0) => Y1_0_port);
   mux010 : MUX21_GENERIC_NBIT16_6 port map( A(15) => Y0_15_port, A(14) => 
                           Y0_14_port, A(13) => Y0_13_port, A(12) => Y0_12_port
                           , A(11) => Y0_11_port, A(10) => Y0_10_port, A(9) => 
                           Y0_9_port, A(8) => Y0_8_port, A(7) => Y0_7_port, 
                           A(6) => Y0_6_port, A(5) => Y0_5_port, A(4) => 
                           Y0_4_port, A(3) => Y0_3_port, A(2) => Y0_2_port, 
                           A(1) => Y0_1_port, A(0) => Y0_0_port, B(15) => 
                           Y1_15_port, B(14) => Y1_14_port, B(13) => Y1_13_port
                           , B(12) => Y1_12_port, B(11) => Y1_11_port, B(10) =>
                           Y1_10_port, B(9) => Y1_9_port, B(8) => Y1_8_port, 
                           B(7) => Y1_7_port, B(6) => Y1_6_port, B(5) => 
                           Y1_5_port, B(4) => Y1_4_port, B(3) => Y1_3_port, 
                           B(2) => Y1_2_port, B(1) => Y1_1_port, B(0) => 
                           Y1_0_port, SEL => SEL(1), Y(15) => Y2_15_port, Y(14)
                           => Y2_14_port, Y(13) => Y2_13_port, Y(12) => 
                           Y2_12_port, Y(11) => Y2_11_port, Y(10) => Y2_10_port
                           , Y(9) => Y2_9_port, Y(8) => Y2_8_port, Y(7) => 
                           Y2_7_port, Y(6) => Y2_6_port, Y(5) => Y2_5_port, 
                           Y(4) => Y2_4_port, Y(3) => Y2_3_port, Y(2) => 
                           Y2_2_port, Y(1) => Y2_1_port, Y(0) => Y2_0_port);
   mux001 : MUX21_GENERIC_NBIT16_5 port map( A(15) => Y2_15_port, A(14) => 
                           Y2_14_port, A(13) => Y2_13_port, A(12) => Y2_12_port
                           , A(11) => Y2_11_port, A(10) => Y2_10_port, A(9) => 
                           Y2_9_port, A(8) => Y2_8_port, A(7) => Y2_7_port, 
                           A(6) => Y2_6_port, A(5) => Y2_5_port, A(4) => 
                           Y2_4_port, A(3) => Y2_3_port, A(2) => Y2_2_port, 
                           A(1) => Y2_1_port, A(0) => Y2_0_port, B(15) => 
                           A4(15), B(14) => A4(14), B(13) => A4(13), B(12) => 
                           A4(12), B(11) => A4(11), B(10) => A4(10), B(9) => 
                           A4(9), B(8) => A4(8), B(7) => A4(7), B(6) => A4(6), 
                           B(5) => A4(5), B(4) => A4(4), B(3) => A4(3), B(2) =>
                           A4(2), B(1) => A4(1), B(0) => A4(0), SEL => SEL(0), 
                           Y(15) => Y(15), Y(14) => Y(14), Y(13) => Y(13), 
                           Y(12) => Y(12), Y(11) => Y(11), Y(10) => Y(10), Y(9)
                           => Y(9), Y(8) => Y(8), Y(7) => Y(7), Y(6) => Y(6), 
                           Y(5) => Y(5), Y(4) => Y(4), Y(3) => Y(3), Y(2) => 
                           Y(2), Y(1) => Y(1), Y(0) => Y(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX51_GENERIC_NBIT16_1 is

   port( A0, A1, A2, A3, A4 : in std_logic_vector (15 downto 0);  SEL : in 
         std_logic_vector (2 downto 0);  Y : out std_logic_vector (15 downto 0)
         );

end MUX51_GENERIC_NBIT16_1;

architecture SYN_STRUCTURAL of MUX51_GENERIC_NBIT16_1 is

   component MUX21_GENERIC_NBIT16_1
      port( A, B : in std_logic_vector (15 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (15 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT16_2
      port( A, B : in std_logic_vector (15 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (15 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT16_3
      port( A, B : in std_logic_vector (15 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (15 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT16_4
      port( A, B : in std_logic_vector (15 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (15 downto 0));
   end component;
   
   signal Y0_15_port, Y0_14_port, Y0_13_port, Y0_12_port, Y0_11_port, 
      Y0_10_port, Y0_9_port, Y0_8_port, Y0_7_port, Y0_6_port, Y0_5_port, 
      Y0_4_port, Y0_3_port, Y0_2_port, Y0_1_port, Y0_0_port, Y1_15_port, 
      Y1_14_port, Y1_13_port, Y1_12_port, Y1_11_port, Y1_10_port, Y1_9_port, 
      Y1_8_port, Y1_7_port, Y1_6_port, Y1_5_port, Y1_4_port, Y1_3_port, 
      Y1_2_port, Y1_1_port, Y1_0_port, Y2_15_port, Y2_14_port, Y2_13_port, 
      Y2_12_port, Y2_11_port, Y2_10_port, Y2_9_port, Y2_8_port, Y2_7_port, 
      Y2_6_port, Y2_5_port, Y2_4_port, Y2_3_port, Y2_2_port, Y2_1_port, 
      Y2_0_port : std_logic;

begin
   
   mux000 : MUX21_GENERIC_NBIT16_4 port map( A(15) => A0(15), A(14) => A0(14), 
                           A(13) => A0(13), A(12) => A0(12), A(11) => A0(11), 
                           A(10) => A0(10), A(9) => A0(9), A(8) => A0(8), A(7) 
                           => A0(7), A(6) => A0(6), A(5) => A0(5), A(4) => 
                           A0(4), A(3) => A0(3), A(2) => A0(2), A(1) => A0(1), 
                           A(0) => A0(0), B(15) => A1(15), B(14) => A1(14), 
                           B(13) => A1(13), B(12) => A1(12), B(11) => A1(11), 
                           B(10) => A1(10), B(9) => A1(9), B(8) => A1(8), B(7) 
                           => A1(7), B(6) => A1(6), B(5) => A1(5), B(4) => 
                           A1(4), B(3) => A1(3), B(2) => A1(2), B(1) => A1(1), 
                           B(0) => A1(0), SEL => SEL(2), Y(15) => Y0_15_port, 
                           Y(14) => Y0_14_port, Y(13) => Y0_13_port, Y(12) => 
                           Y0_12_port, Y(11) => Y0_11_port, Y(10) => Y0_10_port
                           , Y(9) => Y0_9_port, Y(8) => Y0_8_port, Y(7) => 
                           Y0_7_port, Y(6) => Y0_6_port, Y(5) => Y0_5_port, 
                           Y(4) => Y0_4_port, Y(3) => Y0_3_port, Y(2) => 
                           Y0_2_port, Y(1) => Y0_1_port, Y(0) => Y0_0_port);
   mux100 : MUX21_GENERIC_NBIT16_3 port map( A(15) => A2(15), A(14) => A2(14), 
                           A(13) => A2(13), A(12) => A2(12), A(11) => A2(11), 
                           A(10) => A2(10), A(9) => A2(9), A(8) => A2(8), A(7) 
                           => A2(7), A(6) => A2(6), A(5) => A2(5), A(4) => 
                           A2(4), A(3) => A2(3), A(2) => A2(2), A(1) => A2(1), 
                           A(0) => A2(0), B(15) => A3(15), B(14) => A3(14), 
                           B(13) => A3(13), B(12) => A3(12), B(11) => A3(11), 
                           B(10) => A3(10), B(9) => A3(9), B(8) => A3(8), B(7) 
                           => A3(7), B(6) => A3(6), B(5) => A3(5), B(4) => 
                           A3(4), B(3) => A3(3), B(2) => A3(2), B(1) => A3(1), 
                           B(0) => A3(0), SEL => SEL(2), Y(15) => Y1_15_port, 
                           Y(14) => Y1_14_port, Y(13) => Y1_13_port, Y(12) => 
                           Y1_12_port, Y(11) => Y1_11_port, Y(10) => Y1_10_port
                           , Y(9) => Y1_9_port, Y(8) => Y1_8_port, Y(7) => 
                           Y1_7_port, Y(6) => Y1_6_port, Y(5) => Y1_5_port, 
                           Y(4) => Y1_4_port, Y(3) => Y1_3_port, Y(2) => 
                           Y1_2_port, Y(1) => Y1_1_port, Y(0) => Y1_0_port);
   mux010 : MUX21_GENERIC_NBIT16_2 port map( A(15) => Y0_15_port, A(14) => 
                           Y0_14_port, A(13) => Y0_13_port, A(12) => Y0_12_port
                           , A(11) => Y0_11_port, A(10) => Y0_10_port, A(9) => 
                           Y0_9_port, A(8) => Y0_8_port, A(7) => Y0_7_port, 
                           A(6) => Y0_6_port, A(5) => Y0_5_port, A(4) => 
                           Y0_4_port, A(3) => Y0_3_port, A(2) => Y0_2_port, 
                           A(1) => Y0_1_port, A(0) => Y0_0_port, B(15) => 
                           Y1_15_port, B(14) => Y1_14_port, B(13) => Y1_13_port
                           , B(12) => Y1_12_port, B(11) => Y1_11_port, B(10) =>
                           Y1_10_port, B(9) => Y1_9_port, B(8) => Y1_8_port, 
                           B(7) => Y1_7_port, B(6) => Y1_6_port, B(5) => 
                           Y1_5_port, B(4) => Y1_4_port, B(3) => Y1_3_port, 
                           B(2) => Y1_2_port, B(1) => Y1_1_port, B(0) => 
                           Y1_0_port, SEL => SEL(1), Y(15) => Y2_15_port, Y(14)
                           => Y2_14_port, Y(13) => Y2_13_port, Y(12) => 
                           Y2_12_port, Y(11) => Y2_11_port, Y(10) => Y2_10_port
                           , Y(9) => Y2_9_port, Y(8) => Y2_8_port, Y(7) => 
                           Y2_7_port, Y(6) => Y2_6_port, Y(5) => Y2_5_port, 
                           Y(4) => Y2_4_port, Y(3) => Y2_3_port, Y(2) => 
                           Y2_2_port, Y(1) => Y2_1_port, Y(0) => Y2_0_port);
   mux001 : MUX21_GENERIC_NBIT16_1 port map( A(15) => Y2_15_port, A(14) => 
                           Y2_14_port, A(13) => Y2_13_port, A(12) => Y2_12_port
                           , A(11) => Y2_11_port, A(10) => Y2_10_port, A(9) => 
                           Y2_9_port, A(8) => Y2_8_port, A(7) => Y2_7_port, 
                           A(6) => Y2_6_port, A(5) => Y2_5_port, A(4) => 
                           Y2_4_port, A(3) => Y2_3_port, A(2) => Y2_2_port, 
                           A(1) => Y2_1_port, A(0) => Y2_0_port, B(15) => 
                           A4(15), B(14) => A4(14), B(13) => A4(13), B(12) => 
                           A4(12), B(11) => A4(11), B(10) => A4(10), B(9) => 
                           A4(9), B(8) => A4(8), B(7) => A4(7), B(6) => A4(6), 
                           B(5) => A4(5), B(4) => A4(4), B(3) => A4(3), B(2) =>
                           A4(2), B(1) => A4(1), B(0) => A4(0), SEL => SEL(0), 
                           Y(15) => Y(15), Y(14) => Y(14), Y(13) => Y(13), 
                           Y(12) => Y(12), Y(11) => Y(11), Y(10) => Y(10), Y(9)
                           => Y(9), Y(8) => Y(8), Y(7) => Y(7), Y(6) => Y(6), 
                           Y(5) => Y(5), Y(4) => Y(4), Y(3) => Y(3), Y(2) => 
                           Y(2), Y(1) => Y(1), Y(0) => Y(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity SETTLER_NBIT16_3 is

   port( A : in std_logic_vector (15 downto 0);  Y0, Y1, Y2, Y3, Y4, Y5 : out 
         std_logic_vector (15 downto 0));

end SETTLER_NBIT16_3;

architecture SYN_BEHAVIOR of SETTLER_NBIT16_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component SETTLER_NBIT16_3_DW01_inc_0
      port( A : in std_logic_vector (15 downto 0);  SUM : out std_logic_vector 
            (15 downto 0));
   end component;
   
   signal X_Logic0_port, Y2_1_port, Y2_2_port, Y2_3_port, Y2_4_port, Y2_5_port,
      Y2_6_port, Y2_7_port, Y2_8_port, Y2_9_port, Y2_10_port, Y2_11_port, 
      Y2_12_port, Y2_13_port, Y2_14_port, Y2_15_port, n17, n18, n19, n20, n21, 
      n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36
      , n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n_1008 : 
      std_logic;

begin
   Y0 <= ( X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port );
   Y1 <= ( A(15), A(14), A(13), A(12), A(11), A(10), A(9), A(8), A(7), A(6), 
      A(5), A(4), A(3), A(2), A(1), A(0) );
   Y2 <= ( Y2_15_port, Y2_14_port, Y2_13_port, Y2_12_port, Y2_11_port, 
      Y2_10_port, Y2_9_port, Y2_8_port, Y2_7_port, Y2_6_port, Y2_5_port, 
      Y2_4_port, Y2_3_port, Y2_2_port, Y2_1_port, A(0) );
   Y3 <= ( A(14), A(13), A(12), A(11), A(10), A(9), A(8), A(7), A(6), A(5), 
      A(4), A(3), A(2), A(1), A(0), X_Logic0_port );
   Y5 <= ( A(13), A(12), A(11), A(10), A(9), A(8), A(7), A(6), A(5), A(4), A(3)
      , A(2), A(1), A(0), X_Logic0_port, X_Logic0_port );
   
   X_Logic0_port <= '0';
   n47 <= '1';
   add_22 : SETTLER_NBIT16_3_DW01_inc_0 port map( A(15) => n39, A(14) => n40, 
                           A(13) => n41, A(12) => n42, A(11) => n43, A(10) => 
                           n44, A(9) => n37, A(8) => n36, A(7) => n35, A(6) => 
                           n34, A(5) => n33, A(4) => n32, A(3) => n31, A(2) => 
                           n45, A(1) => n46, A(0) => n47, SUM(15) => Y4(15), 
                           SUM(14) => Y4(14), SUM(13) => Y4(13), SUM(12) => 
                           Y4(12), SUM(11) => Y4(11), SUM(10) => Y4(10), SUM(9)
                           => Y4(9), SUM(8) => Y4(8), SUM(7) => Y4(7), SUM(6) 
                           => Y4(6), SUM(5) => Y4(5), SUM(4) => Y4(4), SUM(3) 
                           => Y4(3), SUM(2) => Y4(2), SUM(1) => Y4(1), SUM(0) 
                           => n_1008);
   U3 : XOR2_X1 port map( A => n45, B => n46, Z => Y2_1_port);
   U4 : XOR2_X1 port map( A => n31, B => n29, Z => Y2_2_port);
   U6 : XOR2_X1 port map( A => n32, B => n17, Z => Y2_3_port);
   U7 : XOR2_X1 port map( A => n33, B => n18, Z => Y2_4_port);
   U8 : XOR2_X1 port map( A => n34, B => n19, Z => Y2_5_port);
   U9 : XOR2_X1 port map( A => n35, B => n20, Z => Y2_6_port);
   U10 : XOR2_X1 port map( A => n36, B => n21, Z => Y2_7_port);
   U11 : XOR2_X1 port map( A => n37, B => n22, Z => Y2_8_port);
   U12 : XOR2_X1 port map( A => n44, B => n23, Z => Y2_9_port);
   U13 : XOR2_X1 port map( A => n43, B => n24, Z => Y2_10_port);
   U14 : XOR2_X1 port map( A => n42, B => n25, Z => Y2_11_port);
   U15 : XOR2_X1 port map( A => n41, B => n26, Z => Y2_12_port);
   U16 : XOR2_X1 port map( A => n40, B => n27, Z => Y2_13_port);
   U17 : XOR2_X1 port map( A => n39, B => n28, Z => Y2_14_port);
   U18 : XNOR2_X1 port map( A => n38, B => n30, ZN => Y2_15_port);
   U19 : AND2_X1 port map( A1 => n31, A2 => n29, ZN => n17);
   U20 : AND2_X1 port map( A1 => n32, A2 => n17, ZN => n18);
   U21 : AND2_X1 port map( A1 => n33, A2 => n18, ZN => n19);
   U22 : AND2_X1 port map( A1 => n34, A2 => n19, ZN => n20);
   U23 : AND2_X1 port map( A1 => n35, A2 => n20, ZN => n21);
   U24 : AND2_X1 port map( A1 => n36, A2 => n21, ZN => n22);
   U25 : AND2_X1 port map( A1 => n37, A2 => n22, ZN => n23);
   U26 : AND2_X1 port map( A1 => n44, A2 => n23, ZN => n24);
   U27 : AND2_X1 port map( A1 => n43, A2 => n24, ZN => n25);
   U28 : AND2_X1 port map( A1 => n42, A2 => n25, ZN => n26);
   U29 : AND2_X1 port map( A1 => n41, A2 => n26, ZN => n27);
   U30 : AND2_X1 port map( A1 => n40, A2 => n27, ZN => n28);
   U31 : AND2_X1 port map( A1 => n45, A2 => n46, ZN => n29);
   U32 : NAND2_X1 port map( A1 => n39, A2 => n28, ZN => n30);
   U33 : INV_X1 port map( A => A(15), ZN => n38);
   U34 : INV_X1 port map( A => A(0), ZN => n46);
   U35 : INV_X1 port map( A => A(1), ZN => n45);
   U36 : INV_X1 port map( A => A(9), ZN => n44);
   U37 : INV_X1 port map( A => A(10), ZN => n43);
   U38 : INV_X1 port map( A => A(11), ZN => n42);
   U39 : INV_X1 port map( A => A(12), ZN => n41);
   U40 : INV_X1 port map( A => A(13), ZN => n40);
   U41 : INV_X1 port map( A => A(14), ZN => n39);
   U42 : INV_X1 port map( A => A(8), ZN => n37);
   U43 : INV_X1 port map( A => A(7), ZN => n36);
   U44 : INV_X1 port map( A => A(6), ZN => n35);
   U45 : INV_X1 port map( A => A(5), ZN => n34);
   U46 : INV_X1 port map( A => A(4), ZN => n33);
   U47 : INV_X1 port map( A => A(3), ZN => n32);
   U48 : INV_X1 port map( A => A(2), ZN => n31);
   Y4(0) <= '0';

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity SETTLER_NBIT16_2 is

   port( A : in std_logic_vector (15 downto 0);  Y0, Y1, Y2, Y3, Y4, Y5 : out 
         std_logic_vector (15 downto 0));

end SETTLER_NBIT16_2;

architecture SYN_BEHAVIOR of SETTLER_NBIT16_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component SETTLER_NBIT16_2_DW01_inc_0
      port( A : in std_logic_vector (15 downto 0);  SUM : out std_logic_vector 
            (15 downto 0));
   end component;
   
   signal X_Logic0_port, Y2_1_port, Y2_2_port, Y2_3_port, Y2_4_port, Y2_5_port,
      Y2_6_port, Y2_7_port, Y2_8_port, Y2_9_port, Y2_10_port, Y2_11_port, 
      Y2_12_port, Y2_13_port, Y2_14_port, Y2_15_port, n17, n18, n19, n20, n21, 
      n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36
      , n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n_1009 : 
      std_logic;

begin
   Y0 <= ( X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port );
   Y1 <= ( A(15), A(14), A(13), A(12), A(11), A(10), A(9), A(8), A(7), A(6), 
      A(5), A(4), A(3), A(2), A(1), A(0) );
   Y2 <= ( Y2_15_port, Y2_14_port, Y2_13_port, Y2_12_port, Y2_11_port, 
      Y2_10_port, Y2_9_port, Y2_8_port, Y2_7_port, Y2_6_port, Y2_5_port, 
      Y2_4_port, Y2_3_port, Y2_2_port, Y2_1_port, A(0) );
   Y3 <= ( A(14), A(13), A(12), A(11), A(10), A(9), A(8), A(7), A(6), A(5), 
      A(4), A(3), A(2), A(1), A(0), X_Logic0_port );
   Y5 <= ( A(13), A(12), A(11), A(10), A(9), A(8), A(7), A(6), A(5), A(4), A(3)
      , A(2), A(1), A(0), X_Logic0_port, X_Logic0_port );
   
   X_Logic0_port <= '0';
   n47 <= '1';
   add_22 : SETTLER_NBIT16_2_DW01_inc_0 port map( A(15) => n39, A(14) => n40, 
                           A(13) => n41, A(12) => n42, A(11) => n37, A(10) => 
                           n36, A(9) => n35, A(8) => n34, A(7) => n33, A(6) => 
                           n32, A(5) => n31, A(4) => n43, A(3) => n44, A(2) => 
                           n45, A(1) => n46, A(0) => n47, SUM(15) => Y4(15), 
                           SUM(14) => Y4(14), SUM(13) => Y4(13), SUM(12) => 
                           Y4(12), SUM(11) => Y4(11), SUM(10) => Y4(10), SUM(9)
                           => Y4(9), SUM(8) => Y4(8), SUM(7) => Y4(7), SUM(6) 
                           => Y4(6), SUM(5) => Y4(5), SUM(4) => Y4(4), SUM(3) 
                           => Y4(3), SUM(2) => Y4(2), SUM(1) => Y4(1), SUM(0) 
                           => n_1009);
   U3 : XOR2_X1 port map( A => n45, B => n46, Z => Y2_1_port);
   U4 : XOR2_X1 port map( A => n44, B => n29, Z => Y2_2_port);
   U6 : XOR2_X1 port map( A => n43, B => n28, Z => Y2_3_port);
   U7 : XOR2_X1 port map( A => n31, B => n27, Z => Y2_4_port);
   U8 : XOR2_X1 port map( A => n32, B => n17, Z => Y2_5_port);
   U9 : XOR2_X1 port map( A => n33, B => n18, Z => Y2_6_port);
   U10 : XOR2_X1 port map( A => n34, B => n19, Z => Y2_7_port);
   U11 : XOR2_X1 port map( A => n35, B => n20, Z => Y2_8_port);
   U12 : XOR2_X1 port map( A => n36, B => n21, Z => Y2_9_port);
   U13 : XOR2_X1 port map( A => n37, B => n22, Z => Y2_10_port);
   U14 : XOR2_X1 port map( A => n42, B => n23, Z => Y2_11_port);
   U15 : XOR2_X1 port map( A => n41, B => n24, Z => Y2_12_port);
   U16 : XOR2_X1 port map( A => n40, B => n25, Z => Y2_13_port);
   U17 : XOR2_X1 port map( A => n39, B => n26, Z => Y2_14_port);
   U18 : XNOR2_X1 port map( A => n38, B => n30, ZN => Y2_15_port);
   U19 : AND2_X1 port map( A1 => n31, A2 => n27, ZN => n17);
   U20 : AND2_X1 port map( A1 => n32, A2 => n17, ZN => n18);
   U21 : AND2_X1 port map( A1 => n33, A2 => n18, ZN => n19);
   U22 : AND2_X1 port map( A1 => n34, A2 => n19, ZN => n20);
   U23 : AND2_X1 port map( A1 => n35, A2 => n20, ZN => n21);
   U24 : AND2_X1 port map( A1 => n36, A2 => n21, ZN => n22);
   U25 : AND2_X1 port map( A1 => n37, A2 => n22, ZN => n23);
   U26 : AND2_X1 port map( A1 => n42, A2 => n23, ZN => n24);
   U27 : AND2_X1 port map( A1 => n41, A2 => n24, ZN => n25);
   U28 : AND2_X1 port map( A1 => n40, A2 => n25, ZN => n26);
   U29 : AND2_X1 port map( A1 => n43, A2 => n28, ZN => n27);
   U30 : AND2_X1 port map( A1 => n44, A2 => n29, ZN => n28);
   U31 : AND2_X1 port map( A1 => n45, A2 => n46, ZN => n29);
   U32 : NAND2_X1 port map( A1 => n39, A2 => n26, ZN => n30);
   U33 : INV_X1 port map( A => A(15), ZN => n38);
   U34 : INV_X1 port map( A => A(0), ZN => n46);
   U35 : INV_X1 port map( A => A(1), ZN => n45);
   U36 : INV_X1 port map( A => A(2), ZN => n44);
   U37 : INV_X1 port map( A => A(3), ZN => n43);
   U38 : INV_X1 port map( A => A(11), ZN => n42);
   U39 : INV_X1 port map( A => A(12), ZN => n41);
   U40 : INV_X1 port map( A => A(13), ZN => n40);
   U41 : INV_X1 port map( A => A(14), ZN => n39);
   U42 : INV_X1 port map( A => A(10), ZN => n37);
   U43 : INV_X1 port map( A => A(9), ZN => n36);
   U44 : INV_X1 port map( A => A(8), ZN => n35);
   U45 : INV_X1 port map( A => A(7), ZN => n34);
   U46 : INV_X1 port map( A => A(6), ZN => n33);
   U47 : INV_X1 port map( A => A(5), ZN => n32);
   U48 : INV_X1 port map( A => A(4), ZN => n31);
   Y4(0) <= '0';

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity SETTLER_NBIT16_1 is

   port( A : in std_logic_vector (15 downto 0);  Y0, Y1, Y2, Y3, Y4, Y5 : out 
         std_logic_vector (15 downto 0));

end SETTLER_NBIT16_1;

architecture SYN_BEHAVIOR of SETTLER_NBIT16_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component SETTLER_NBIT16_1_DW01_inc_0
      port( A : in std_logic_vector (15 downto 0);  SUM : out std_logic_vector 
            (15 downto 0));
   end component;
   
   signal X_Logic0_port, Y2_1_port, Y2_2_port, Y2_3_port, Y2_4_port, Y2_5_port,
      Y2_6_port, Y2_7_port, Y2_8_port, Y2_9_port, Y2_10_port, Y2_11_port, 
      Y2_12_port, Y2_13_port, Y2_14_port, Y2_15_port, n17, n18, n19, n20, n21, 
      n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36
      , n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n_1010 : 
      std_logic;

begin
   Y0 <= ( X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port );
   Y1 <= ( A(15), A(14), A(13), A(12), A(11), A(10), A(9), A(8), A(7), A(6), 
      A(5), A(4), A(3), A(2), A(1), A(0) );
   Y2 <= ( Y2_15_port, Y2_14_port, Y2_13_port, Y2_12_port, Y2_11_port, 
      Y2_10_port, Y2_9_port, Y2_8_port, Y2_7_port, Y2_6_port, Y2_5_port, 
      Y2_4_port, Y2_3_port, Y2_2_port, Y2_1_port, A(0) );
   Y3 <= ( A(14), A(13), A(12), A(11), A(10), A(9), A(8), A(7), A(6), A(5), 
      A(4), A(3), A(2), A(1), A(0), X_Logic0_port );
   Y5 <= ( A(13), A(12), A(11), A(10), A(9), A(8), A(7), A(6), A(5), A(4), A(3)
      , A(2), A(1), A(0), X_Logic0_port, X_Logic0_port );
   
   X_Logic0_port <= '0';
   n47 <= '1';
   add_22 : SETTLER_NBIT16_1_DW01_inc_0 port map( A(15) => n39, A(14) => n40, 
                           A(13) => n37, A(12) => n36, A(11) => n35, A(10) => 
                           n34, A(9) => n33, A(8) => n32, A(7) => n31, A(6) => 
                           n41, A(5) => n42, A(4) => n45, A(3) => n46, A(2) => 
                           n43, A(1) => n44, A(0) => n47, SUM(15) => Y4(15), 
                           SUM(14) => Y4(14), SUM(13) => Y4(13), SUM(12) => 
                           Y4(12), SUM(11) => Y4(11), SUM(10) => Y4(10), SUM(9)
                           => Y4(9), SUM(8) => Y4(8), SUM(7) => Y4(7), SUM(6) 
                           => Y4(6), SUM(5) => Y4(5), SUM(4) => Y4(4), SUM(3) 
                           => Y4(3), SUM(2) => Y4(2), SUM(1) => Y4(1), SUM(0) 
                           => n_1010);
   U3 : XOR2_X1 port map( A => n43, B => n44, Z => Y2_1_port);
   U4 : XOR2_X1 port map( A => n46, B => n29, Z => Y2_2_port);
   U6 : XOR2_X1 port map( A => n45, B => n28, Z => Y2_3_port);
   U7 : XOR2_X1 port map( A => n42, B => n25, Z => Y2_4_port);
   U8 : XOR2_X1 port map( A => n41, B => n26, Z => Y2_5_port);
   U9 : XOR2_X1 port map( A => n31, B => n27, Z => Y2_6_port);
   U10 : XOR2_X1 port map( A => n32, B => n17, Z => Y2_7_port);
   U11 : XOR2_X1 port map( A => n33, B => n18, Z => Y2_8_port);
   U12 : XOR2_X1 port map( A => n34, B => n19, Z => Y2_9_port);
   U13 : XOR2_X1 port map( A => n35, B => n20, Z => Y2_10_port);
   U14 : XOR2_X1 port map( A => n36, B => n21, Z => Y2_11_port);
   U15 : XOR2_X1 port map( A => n37, B => n22, Z => Y2_12_port);
   U16 : XOR2_X1 port map( A => n40, B => n23, Z => Y2_13_port);
   U17 : XOR2_X1 port map( A => n39, B => n24, Z => Y2_14_port);
   U18 : XNOR2_X1 port map( A => n38, B => n30, ZN => Y2_15_port);
   U19 : AND2_X1 port map( A1 => n31, A2 => n27, ZN => n17);
   U20 : AND2_X1 port map( A1 => n32, A2 => n17, ZN => n18);
   U21 : AND2_X1 port map( A1 => n33, A2 => n18, ZN => n19);
   U22 : AND2_X1 port map( A1 => n34, A2 => n19, ZN => n20);
   U23 : AND2_X1 port map( A1 => n35, A2 => n20, ZN => n21);
   U24 : AND2_X1 port map( A1 => n36, A2 => n21, ZN => n22);
   U25 : AND2_X1 port map( A1 => n37, A2 => n22, ZN => n23);
   U26 : AND2_X1 port map( A1 => n40, A2 => n23, ZN => n24);
   U27 : AND2_X1 port map( A1 => n45, A2 => n28, ZN => n25);
   U28 : AND2_X1 port map( A1 => n42, A2 => n25, ZN => n26);
   U29 : AND2_X1 port map( A1 => n41, A2 => n26, ZN => n27);
   U30 : AND2_X1 port map( A1 => n46, A2 => n29, ZN => n28);
   U31 : AND2_X1 port map( A1 => n43, A2 => n44, ZN => n29);
   U32 : NAND2_X1 port map( A1 => n39, A2 => n24, ZN => n30);
   U33 : INV_X1 port map( A => A(15), ZN => n38);
   U34 : INV_X1 port map( A => A(2), ZN => n46);
   U35 : INV_X1 port map( A => A(3), ZN => n45);
   U36 : INV_X1 port map( A => A(0), ZN => n44);
   U37 : INV_X1 port map( A => A(1), ZN => n43);
   U38 : INV_X1 port map( A => A(4), ZN => n42);
   U39 : INV_X1 port map( A => A(5), ZN => n41);
   U40 : INV_X1 port map( A => A(13), ZN => n40);
   U41 : INV_X1 port map( A => A(14), ZN => n39);
   U42 : INV_X1 port map( A => A(12), ZN => n37);
   U43 : INV_X1 port map( A => A(11), ZN => n36);
   U44 : INV_X1 port map( A => A(10), ZN => n35);
   U45 : INV_X1 port map( A => A(9), ZN => n34);
   U46 : INV_X1 port map( A => A(8), ZN => n33);
   U47 : INV_X1 port map( A => A(7), ZN => n32);
   U48 : INV_X1 port map( A => A(6), ZN => n31);
   Y4(0) <= '0';

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ENC3TO3_3 is

   port( X : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (2 
         downto 0));

end ENC3TO3_3;

architecture SYN_BEHAVIOR of ENC3TO3_3 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X2
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : MUX2_X2 port map( A => n2, B => n3, S => X(2), Z => Y(1));
   U2 : NAND3_X2 port map( A1 => n3, A2 => n2, A3 => X(2), ZN => Y(0));
   U3 : INV_X4 port map( A => n1, ZN => Y(2));
   U4 : AOI21_X1 port map( B1 => n2, B2 => n3, A => X(2), ZN => n1);
   U5 : NAND2_X1 port map( A1 => X(1), A2 => X(0), ZN => n2);
   U6 : XNOR2_X1 port map( A => X(0), B => X(1), ZN => n3);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ENC3TO3_2 is

   port( X : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (2 
         downto 0));

end ENC3TO3_2;

architecture SYN_BEHAVIOR of ENC3TO3_2 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X2
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : MUX2_X2 port map( A => n2, B => n3, S => X(2), Z => Y(1));
   U2 : NAND3_X2 port map( A1 => n3, A2 => n2, A3 => X(2), ZN => Y(0));
   U3 : INV_X4 port map( A => n1, ZN => Y(2));
   U4 : AOI21_X1 port map( B1 => n2, B2 => n3, A => X(2), ZN => n1);
   U5 : NAND2_X1 port map( A1 => X(1), A2 => X(0), ZN => n2);
   U6 : XNOR2_X1 port map( A => X(0), B => X(1), ZN => n3);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ENC3TO3_1 is

   port( X : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (2 
         downto 0));

end ENC3TO3_1;

architecture SYN_BEHAVIOR of ENC3TO3_1 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X2
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : MUX2_X2 port map( A => n2, B => n3, S => X(2), Z => Y(1));
   U2 : NAND3_X2 port map( A1 => n3, A2 => n2, A3 => X(2), ZN => Y(0));
   U3 : INV_X4 port map( A => n1, ZN => Y(2));
   U4 : AOI21_X1 port map( B1 => n2, B2 => n3, A => X(2), ZN => n1);
   U5 : NAND2_X1 port map( A1 => X(1), A2 => X(0), ZN => n2);
   U6 : XNOR2_X1 port map( A => X(0), B => X(1), ZN => n3);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ND2_0 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_0;

architecture SYN_ARCH2 of ND2_0 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity IV_0 is

   port( A : in std_logic;  Y : out std_logic);

end IV_0;

architecture SYN_BEHAVIORAL of IV_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_0 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_0;

architecture SYN_STRUCTURAL of MUX21_0 is

   component ND2_766
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_767
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_0
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_0
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_0 port map( A => S, Y => SB);
   UND1 : ND2_0 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_767 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_766 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity FA_0 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_0;

architecture SYN_Behavioural of FA_0 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => c_in, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => c_out);
   U3 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n1, B2 => c_in, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n1);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX21_GENERIC_NBIT16_0 is

   port( A, B : in std_logic_vector (15 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (15 downto 0));

end MUX21_GENERIC_NBIT16_0;

architecture SYN_STRUCTURAL of MUX21_GENERIC_NBIT16_0 is

   component MUX21_241
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_242
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_243
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_244
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_245
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_246
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_247
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_248
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_249
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_250
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_251
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_252
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_253
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_254
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_255
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_0
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUX21GENI_0 : MUX21_0 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUX21GENI_1 : MUX21_255 port map( A => A(1), B => B(1), S => SEL, Y => Y(1))
                           ;
   MUX21GENI_2 : MUX21_254 port map( A => A(2), B => B(2), S => SEL, Y => Y(2))
                           ;
   MUX21GENI_3 : MUX21_253 port map( A => A(3), B => B(3), S => SEL, Y => Y(3))
                           ;
   MUX21GENI_4 : MUX21_252 port map( A => A(4), B => B(4), S => SEL, Y => Y(4))
                           ;
   MUX21GENI_5 : MUX21_251 port map( A => A(5), B => B(5), S => SEL, Y => Y(5))
                           ;
   MUX21GENI_6 : MUX21_250 port map( A => A(6), B => B(6), S => SEL, Y => Y(6))
                           ;
   MUX21GENI_7 : MUX21_249 port map( A => A(7), B => B(7), S => SEL, Y => Y(7))
                           ;
   MUX21GENI_8 : MUX21_248 port map( A => A(8), B => B(8), S => SEL, Y => Y(8))
                           ;
   MUX21GENI_9 : MUX21_247 port map( A => A(9), B => B(9), S => SEL, Y => Y(9))
                           ;
   MUX21GENI_10 : MUX21_246 port map( A => A(10), B => B(10), S => SEL, Y => 
                           Y(10));
   MUX21GENI_11 : MUX21_245 port map( A => A(11), B => B(11), S => SEL, Y => 
                           Y(11));
   MUX21GENI_12 : MUX21_244 port map( A => A(12), B => B(12), S => SEL, Y => 
                           Y(12));
   MUX21GENI_13 : MUX21_243 port map( A => A(13), B => B(13), S => SEL, Y => 
                           Y(13));
   MUX21GENI_14 : MUX21_242 port map( A => A(14), B => B(14), S => SEL, Y => 
                           Y(14));
   MUX21GENI_15 : MUX21_241 port map( A => A(15), B => B(15), S => SEL, Y => 
                           Y(15));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity RCA_size16_0 is

   port( a, b : in std_logic_vector (15 downto 0);  c_in : in std_logic;  c_out
         : out std_logic;  sum : out std_logic_vector (15 downto 0));

end RCA_size16_0;

architecture SYN_Structural of RCA_size16_0 is

   component FA_33
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_34
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_35
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_36
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_37
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_38
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_39
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_40
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_41
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_42
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_43
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_44
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_45
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_46
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_47
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_0
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   signal temp_15_port, temp_14_port, temp_13_port, temp_12_port, temp_11_port,
      temp_10_port, temp_9_port, temp_8_port, temp_7_port, temp_6_port, 
      temp_5_port, temp_4_port, temp_3_port, temp_2_port, temp_1_port : 
      std_logic;

begin
   
   fa_i_0 : FA_0 port map( a => a(0), b => b(0), c_in => c_in, c_out => 
                           temp_1_port, s => sum(0));
   fa_i_1 : FA_47 port map( a => a(1), b => b(1), c_in => temp_1_port, c_out =>
                           temp_2_port, s => sum(1));
   fa_i_2 : FA_46 port map( a => a(2), b => b(2), c_in => temp_2_port, c_out =>
                           temp_3_port, s => sum(2));
   fa_i_3 : FA_45 port map( a => a(3), b => b(3), c_in => temp_3_port, c_out =>
                           temp_4_port, s => sum(3));
   fa_i_4 : FA_44 port map( a => a(4), b => b(4), c_in => temp_4_port, c_out =>
                           temp_5_port, s => sum(4));
   fa_i_5 : FA_43 port map( a => a(5), b => b(5), c_in => temp_5_port, c_out =>
                           temp_6_port, s => sum(5));
   fa_i_6 : FA_42 port map( a => a(6), b => b(6), c_in => temp_6_port, c_out =>
                           temp_7_port, s => sum(6));
   fa_i_7 : FA_41 port map( a => a(7), b => b(7), c_in => temp_7_port, c_out =>
                           temp_8_port, s => sum(7));
   fa_i_8 : FA_40 port map( a => a(8), b => b(8), c_in => temp_8_port, c_out =>
                           temp_9_port, s => sum(8));
   fa_i_9 : FA_39 port map( a => a(9), b => b(9), c_in => temp_9_port, c_out =>
                           temp_10_port, s => sum(9));
   fa_i_10 : FA_38 port map( a => a(10), b => b(10), c_in => temp_10_port, 
                           c_out => temp_11_port, s => sum(10));
   fa_i_11 : FA_37 port map( a => a(11), b => b(11), c_in => temp_11_port, 
                           c_out => temp_12_port, s => sum(11));
   fa_i_12 : FA_36 port map( a => a(12), b => b(12), c_in => temp_12_port, 
                           c_out => temp_13_port, s => sum(12));
   fa_i_13 : FA_35 port map( a => a(13), b => b(13), c_in => temp_13_port, 
                           c_out => temp_14_port, s => sum(13));
   fa_i_14 : FA_34 port map( a => a(14), b => b(14), c_in => temp_14_port, 
                           c_out => temp_15_port, s => sum(14));
   fa_i_15 : FA_33 port map( a => a(15), b => b(15), c_in => temp_15_port, 
                           c_out => c_out, s => sum(15));

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity MUX51_GENERIC_NBIT16_0 is

   port( A0, A1, A2, A3, A4 : in std_logic_vector (15 downto 0);  SEL : in 
         std_logic_vector (2 downto 0);  Y : out std_logic_vector (15 downto 0)
         );

end MUX51_GENERIC_NBIT16_0;

architecture SYN_STRUCTURAL of MUX51_GENERIC_NBIT16_0 is

   component MUX21_GENERIC_NBIT16_13
      port( A, B : in std_logic_vector (15 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (15 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT16_14
      port( A, B : in std_logic_vector (15 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (15 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT16_15
      port( A, B : in std_logic_vector (15 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (15 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT16_0
      port( A, B : in std_logic_vector (15 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (15 downto 0));
   end component;
   
   signal Y0_15_port, Y0_14_port, Y0_13_port, Y0_12_port, Y0_11_port, 
      Y0_10_port, Y0_9_port, Y0_8_port, Y0_7_port, Y0_6_port, Y0_5_port, 
      Y0_4_port, Y0_3_port, Y0_2_port, Y0_1_port, Y0_0_port, Y1_15_port, 
      Y1_14_port, Y1_13_port, Y1_12_port, Y1_11_port, Y1_10_port, Y1_9_port, 
      Y1_8_port, Y1_7_port, Y1_6_port, Y1_5_port, Y1_4_port, Y1_3_port, 
      Y1_2_port, Y1_1_port, Y1_0_port, Y2_15_port, Y2_14_port, Y2_13_port, 
      Y2_12_port, Y2_11_port, Y2_10_port, Y2_9_port, Y2_8_port, Y2_7_port, 
      Y2_6_port, Y2_5_port, Y2_4_port, Y2_3_port, Y2_2_port, Y2_1_port, 
      Y2_0_port : std_logic;

begin
   
   mux000 : MUX21_GENERIC_NBIT16_0 port map( A(15) => A0(15), A(14) => A0(14), 
                           A(13) => A0(13), A(12) => A0(12), A(11) => A0(11), 
                           A(10) => A0(10), A(9) => A0(9), A(8) => A0(8), A(7) 
                           => A0(7), A(6) => A0(6), A(5) => A0(5), A(4) => 
                           A0(4), A(3) => A0(3), A(2) => A0(2), A(1) => A0(1), 
                           A(0) => A0(0), B(15) => A1(15), B(14) => A1(14), 
                           B(13) => A1(13), B(12) => A1(12), B(11) => A1(11), 
                           B(10) => A1(10), B(9) => A1(9), B(8) => A1(8), B(7) 
                           => A1(7), B(6) => A1(6), B(5) => A1(5), B(4) => 
                           A1(4), B(3) => A1(3), B(2) => A1(2), B(1) => A1(1), 
                           B(0) => A1(0), SEL => SEL(2), Y(15) => Y0_15_port, 
                           Y(14) => Y0_14_port, Y(13) => Y0_13_port, Y(12) => 
                           Y0_12_port, Y(11) => Y0_11_port, Y(10) => Y0_10_port
                           , Y(9) => Y0_9_port, Y(8) => Y0_8_port, Y(7) => 
                           Y0_7_port, Y(6) => Y0_6_port, Y(5) => Y0_5_port, 
                           Y(4) => Y0_4_port, Y(3) => Y0_3_port, Y(2) => 
                           Y0_2_port, Y(1) => Y0_1_port, Y(0) => Y0_0_port);
   mux100 : MUX21_GENERIC_NBIT16_15 port map( A(15) => A2(15), A(14) => A2(14),
                           A(13) => A2(13), A(12) => A2(12), A(11) => A2(11), 
                           A(10) => A2(10), A(9) => A2(9), A(8) => A2(8), A(7) 
                           => A2(7), A(6) => A2(6), A(5) => A2(5), A(4) => 
                           A2(4), A(3) => A2(3), A(2) => A2(2), A(1) => A2(1), 
                           A(0) => A2(0), B(15) => A3(15), B(14) => A3(14), 
                           B(13) => A3(13), B(12) => A3(12), B(11) => A3(11), 
                           B(10) => A3(10), B(9) => A3(9), B(8) => A3(8), B(7) 
                           => A3(7), B(6) => A3(6), B(5) => A3(5), B(4) => 
                           A3(4), B(3) => A3(3), B(2) => A3(2), B(1) => A3(1), 
                           B(0) => A3(0), SEL => SEL(2), Y(15) => Y1_15_port, 
                           Y(14) => Y1_14_port, Y(13) => Y1_13_port, Y(12) => 
                           Y1_12_port, Y(11) => Y1_11_port, Y(10) => Y1_10_port
                           , Y(9) => Y1_9_port, Y(8) => Y1_8_port, Y(7) => 
                           Y1_7_port, Y(6) => Y1_6_port, Y(5) => Y1_5_port, 
                           Y(4) => Y1_4_port, Y(3) => Y1_3_port, Y(2) => 
                           Y1_2_port, Y(1) => Y1_1_port, Y(0) => Y1_0_port);
   mux010 : MUX21_GENERIC_NBIT16_14 port map( A(15) => Y0_15_port, A(14) => 
                           Y0_14_port, A(13) => Y0_13_port, A(12) => Y0_12_port
                           , A(11) => Y0_11_port, A(10) => Y0_10_port, A(9) => 
                           Y0_9_port, A(8) => Y0_8_port, A(7) => Y0_7_port, 
                           A(6) => Y0_6_port, A(5) => Y0_5_port, A(4) => 
                           Y0_4_port, A(3) => Y0_3_port, A(2) => Y0_2_port, 
                           A(1) => Y0_1_port, A(0) => Y0_0_port, B(15) => 
                           Y1_15_port, B(14) => Y1_14_port, B(13) => Y1_13_port
                           , B(12) => Y1_12_port, B(11) => Y1_11_port, B(10) =>
                           Y1_10_port, B(9) => Y1_9_port, B(8) => Y1_8_port, 
                           B(7) => Y1_7_port, B(6) => Y1_6_port, B(5) => 
                           Y1_5_port, B(4) => Y1_4_port, B(3) => Y1_3_port, 
                           B(2) => Y1_2_port, B(1) => Y1_1_port, B(0) => 
                           Y1_0_port, SEL => SEL(1), Y(15) => Y2_15_port, Y(14)
                           => Y2_14_port, Y(13) => Y2_13_port, Y(12) => 
                           Y2_12_port, Y(11) => Y2_11_port, Y(10) => Y2_10_port
                           , Y(9) => Y2_9_port, Y(8) => Y2_8_port, Y(7) => 
                           Y2_7_port, Y(6) => Y2_6_port, Y(5) => Y2_5_port, 
                           Y(4) => Y2_4_port, Y(3) => Y2_3_port, Y(2) => 
                           Y2_2_port, Y(1) => Y2_1_port, Y(0) => Y2_0_port);
   mux001 : MUX21_GENERIC_NBIT16_13 port map( A(15) => Y2_15_port, A(14) => 
                           Y2_14_port, A(13) => Y2_13_port, A(12) => Y2_12_port
                           , A(11) => Y2_11_port, A(10) => Y2_10_port, A(9) => 
                           Y2_9_port, A(8) => Y2_8_port, A(7) => Y2_7_port, 
                           A(6) => Y2_6_port, A(5) => Y2_5_port, A(4) => 
                           Y2_4_port, A(3) => Y2_3_port, A(2) => Y2_2_port, 
                           A(1) => Y2_1_port, A(0) => Y2_0_port, B(15) => 
                           A4(15), B(14) => A4(14), B(13) => A4(13), B(12) => 
                           A4(12), B(11) => A4(11), B(10) => A4(10), B(9) => 
                           A4(9), B(8) => A4(8), B(7) => A4(7), B(6) => A4(6), 
                           B(5) => A4(5), B(4) => A4(4), B(3) => A4(3), B(2) =>
                           A4(2), B(1) => A4(1), B(0) => A4(0), SEL => SEL(0), 
                           Y(15) => Y(15), Y(14) => Y(14), Y(13) => Y(13), 
                           Y(12) => Y(12), Y(11) => Y(11), Y(10) => Y(10), Y(9)
                           => Y(9), Y(8) => Y(8), Y(7) => Y(7), Y(6) => Y(6), 
                           Y(5) => Y(5), Y(4) => Y(4), Y(3) => Y(3), Y(2) => 
                           Y(2), Y(1) => Y(1), Y(0) => Y(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity SETTLER_NBIT16_0 is

   port( A : in std_logic_vector (15 downto 0);  Y0, Y1, Y2, Y3, Y4, Y5 : out 
         std_logic_vector (15 downto 0));

end SETTLER_NBIT16_0;

architecture SYN_BEHAVIOR of SETTLER_NBIT16_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component SETTLER_NBIT16_0_DW01_inc_0
      port( A : in std_logic_vector (15 downto 0);  SUM : out std_logic_vector 
            (15 downto 0));
   end component;
   
   signal X_Logic0_port, n3, Y2_1_port, Y2_2_port, Y2_3_port, Y2_4_port, 
      Y2_5_port, Y2_6_port, Y2_7_port, Y2_8_port, Y2_9_port, Y2_10_port, 
      Y2_11_port, Y2_12_port, Y2_13_port, Y2_14_port, Y2_15_port, n17, n18, n19
      , n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, 
      n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n_1011 :
      std_logic;

begin
   Y0 <= ( X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port );
   Y1 <= ( A(15), A(14), A(13), A(12), A(11), A(10), A(9), A(8), A(7), A(6), 
      A(5), A(4), A(3), A(2), A(1), A(0) );
   Y2 <= ( Y2_15_port, Y2_14_port, Y2_13_port, Y2_12_port, Y2_11_port, 
      Y2_10_port, Y2_9_port, Y2_8_port, Y2_7_port, Y2_6_port, Y2_5_port, 
      Y2_4_port, Y2_3_port, Y2_2_port, Y2_1_port, A(0) );
   Y3 <= ( A(14), A(13), A(12), A(11), A(10), A(9), A(8), A(7), A(6), A(5), 
      A(4), A(3), A(2), A(1), A(0), X_Logic0_port );
   Y5 <= ( A(13), A(12), A(11), A(10), A(9), A(8), A(7), A(6), A(5), A(4), A(3)
      , A(2), A(1), A(0), X_Logic0_port, X_Logic0_port );
   
   X_Logic0_port <= '0';
   n3 <= '1';
   add_22 : SETTLER_NBIT16_0_DW01_inc_0 port map( A(15) => n39, A(14) => n40, 
                           A(13) => n41, A(12) => n42, A(11) => n43, A(10) => 
                           n44, A(9) => n45, A(8) => n46, A(7) => n37, A(6) => 
                           n36, A(5) => n35, A(4) => n34, A(3) => n33, A(2) => 
                           n32, A(1) => n31, A(0) => n3, SUM(15) => Y4(15), 
                           SUM(14) => Y4(14), SUM(13) => Y4(13), SUM(12) => 
                           Y4(12), SUM(11) => Y4(11), SUM(10) => Y4(10), SUM(9)
                           => Y4(9), SUM(8) => Y4(8), SUM(7) => Y4(7), SUM(6) 
                           => Y4(6), SUM(5) => Y4(5), SUM(4) => Y4(4), SUM(3) 
                           => Y4(3), SUM(2) => Y4(2), SUM(1) => Y4(1), SUM(0) 
                           => n_1011);
   U3 : XOR2_X1 port map( A => n32, B => n31, Z => Y2_1_port);
   U4 : XOR2_X1 port map( A => n33, B => n17, Z => Y2_2_port);
   U6 : XOR2_X1 port map( A => n34, B => n18, Z => Y2_3_port);
   U7 : XOR2_X1 port map( A => n35, B => n19, Z => Y2_4_port);
   U8 : XOR2_X1 port map( A => n36, B => n20, Z => Y2_5_port);
   U9 : XOR2_X1 port map( A => n37, B => n21, Z => Y2_6_port);
   U10 : XOR2_X1 port map( A => n46, B => n22, Z => Y2_7_port);
   U11 : XOR2_X1 port map( A => n45, B => n23, Z => Y2_8_port);
   U12 : XOR2_X1 port map( A => n44, B => n24, Z => Y2_9_port);
   U13 : XOR2_X1 port map( A => n43, B => n25, Z => Y2_10_port);
   U14 : XOR2_X1 port map( A => n42, B => n26, Z => Y2_11_port);
   U15 : XOR2_X1 port map( A => n41, B => n27, Z => Y2_12_port);
   U16 : XOR2_X1 port map( A => n40, B => n28, Z => Y2_13_port);
   U17 : XOR2_X1 port map( A => n39, B => n29, Z => Y2_14_port);
   U18 : XNOR2_X1 port map( A => n38, B => n30, ZN => Y2_15_port);
   U19 : AND2_X1 port map( A1 => n32, A2 => n31, ZN => n17);
   U20 : AND2_X1 port map( A1 => n33, A2 => n17, ZN => n18);
   U21 : AND2_X1 port map( A1 => n34, A2 => n18, ZN => n19);
   U22 : AND2_X1 port map( A1 => n35, A2 => n19, ZN => n20);
   U23 : AND2_X1 port map( A1 => n36, A2 => n20, ZN => n21);
   U24 : AND2_X1 port map( A1 => n37, A2 => n21, ZN => n22);
   U25 : AND2_X1 port map( A1 => n46, A2 => n22, ZN => n23);
   U26 : AND2_X1 port map( A1 => n45, A2 => n23, ZN => n24);
   U27 : AND2_X1 port map( A1 => n44, A2 => n24, ZN => n25);
   U28 : AND2_X1 port map( A1 => n43, A2 => n25, ZN => n26);
   U29 : AND2_X1 port map( A1 => n42, A2 => n26, ZN => n27);
   U30 : AND2_X1 port map( A1 => n41, A2 => n27, ZN => n28);
   U31 : AND2_X1 port map( A1 => n40, A2 => n28, ZN => n29);
   U32 : NAND2_X1 port map( A1 => n39, A2 => n29, ZN => n30);
   U33 : INV_X1 port map( A => A(15), ZN => n38);
   U34 : INV_X1 port map( A => A(7), ZN => n46);
   U35 : INV_X1 port map( A => A(8), ZN => n45);
   U36 : INV_X1 port map( A => A(9), ZN => n44);
   U37 : INV_X1 port map( A => A(10), ZN => n43);
   U38 : INV_X1 port map( A => A(11), ZN => n42);
   U39 : INV_X1 port map( A => A(12), ZN => n41);
   U40 : INV_X1 port map( A => A(13), ZN => n40);
   U41 : INV_X1 port map( A => A(14), ZN => n39);
   U42 : INV_X1 port map( A => A(6), ZN => n37);
   U43 : INV_X1 port map( A => A(5), ZN => n36);
   U44 : INV_X1 port map( A => A(4), ZN => n35);
   U45 : INV_X1 port map( A => A(3), ZN => n34);
   U46 : INV_X1 port map( A => A(2), ZN => n33);
   U47 : INV_X1 port map( A => A(1), ZN => n32);
   U48 : INV_X1 port map( A => A(0), ZN => n31);
   Y4(0) <= '0';

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity ENC3TO3_0 is

   port( X : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (2 
         downto 0));

end ENC3TO3_0;

architecture SYN_BEHAVIOR of ENC3TO3_0 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X2
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : MUX2_X2 port map( A => n2, B => n3, S => X(2), Z => Y(1));
   U2 : NAND3_X2 port map( A1 => n3, A2 => n2, A3 => X(2), ZN => Y(0));
   U3 : INV_X4 port map( A => n1, ZN => Y(2));
   U4 : AOI21_X1 port map( B1 => n2, B2 => n3, A => X(2), ZN => n1);
   U5 : NAND2_X1 port map( A1 => X(1), A2 => X(0), ZN => n2);
   U6 : XNOR2_X1 port map( A => X(0), B => X(1), ZN => n3);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT8.all;

entity BOOTHMUL_NBIT8 is

   port( A_mp, B_mp : in std_logic_vector (7 downto 0);  Y_mp : out 
         std_logic_vector (15 downto 0));

end BOOTHMUL_NBIT8;

architecture SYN_STRUCTURAL of BOOTHMUL_NBIT8 is

   component RCA_size16_1
      port( a, b : in std_logic_vector (15 downto 0);  c_in : in std_logic;  
            c_out : out std_logic;  sum : out std_logic_vector (15 downto 0));
   end component;
   
   component MUX51_GENERIC_NBIT16_1
      port( A0, A1, A2, A3, A4 : in std_logic_vector (15 downto 0);  SEL : in 
            std_logic_vector (2 downto 0);  Y : out std_logic_vector (15 downto
            0));
   end component;
   
   component SETTLER_NBIT16_1
      port( A : in std_logic_vector (15 downto 0);  Y0, Y1, Y2, Y3, Y4, Y5 : 
            out std_logic_vector (15 downto 0));
   end component;
   
   component ENC3TO3_1
      port( X : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (2 
            downto 0));
   end component;
   
   component RCA_size16_2
      port( a, b : in std_logic_vector (15 downto 0);  c_in : in std_logic;  
            c_out : out std_logic;  sum : out std_logic_vector (15 downto 0));
   end component;
   
   component MUX51_GENERIC_NBIT16_2
      port( A0, A1, A2, A3, A4 : in std_logic_vector (15 downto 0);  SEL : in 
            std_logic_vector (2 downto 0);  Y : out std_logic_vector (15 downto
            0));
   end component;
   
   component SETTLER_NBIT16_2
      port( A : in std_logic_vector (15 downto 0);  Y0, Y1, Y2, Y3, Y4, Y5 : 
            out std_logic_vector (15 downto 0));
   end component;
   
   component ENC3TO3_2
      port( X : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (2 
            downto 0));
   end component;
   
   component RCA_size16_0
      port( a, b : in std_logic_vector (15 downto 0);  c_in : in std_logic;  
            c_out : out std_logic;  sum : out std_logic_vector (15 downto 0));
   end component;
   
   component MUX51_GENERIC_NBIT16_3
      port( A0, A1, A2, A3, A4 : in std_logic_vector (15 downto 0);  SEL : in 
            std_logic_vector (2 downto 0);  Y : out std_logic_vector (15 downto
            0));
   end component;
   
   component SETTLER_NBIT16_3
      port( A : in std_logic_vector (15 downto 0);  Y0, Y1, Y2, Y3, Y4, Y5 : 
            out std_logic_vector (15 downto 0));
   end component;
   
   component ENC3TO3_3
      port( X : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (2 
            downto 0));
   end component;
   
   component MUX51_GENERIC_NBIT16_0
      port( A0, A1, A2, A3, A4 : in std_logic_vector (15 downto 0);  SEL : in 
            std_logic_vector (2 downto 0);  Y : out std_logic_vector (15 downto
            0));
   end component;
   
   component SETTLER_NBIT16_0
      port( A : in std_logic_vector (15 downto 0);  Y0, Y1, Y2, Y3, Y4, Y5 : 
            out std_logic_vector (15 downto 0));
   end component;
   
   component ENC3TO3_0
      port( X : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (2 
            downto 0));
   end component;
   
   signal X_Logic0_port, set_signal_0_1_15_port, set_signal_0_1_14_port, 
      set_signal_0_1_13_port, set_signal_0_1_12_port, set_signal_0_1_11_port, 
      set_signal_0_1_10_port, set_signal_0_1_9_port, set_signal_0_1_8_port, 
      set_signal_0_1_7_port, set_signal_0_1_6_port, set_signal_0_1_5_port, 
      set_signal_0_1_4_port, set_signal_0_1_3_port, set_signal_0_1_2_port, 
      set_signal_0_1_1_port, set_signal_0_1_0_port, set_signal_0_2_15_port, 
      set_signal_0_2_14_port, set_signal_0_2_13_port, set_signal_0_2_12_port, 
      set_signal_0_2_11_port, set_signal_0_2_10_port, set_signal_0_2_9_port, 
      set_signal_0_2_8_port, set_signal_0_2_7_port, set_signal_0_2_6_port, 
      set_signal_0_2_5_port, set_signal_0_2_4_port, set_signal_0_2_3_port, 
      set_signal_0_2_2_port, set_signal_0_2_1_port, set_signal_0_2_0_port, 
      set_signal_0_3_15_port, set_signal_0_3_14_port, set_signal_0_3_13_port, 
      set_signal_0_3_12_port, set_signal_0_3_11_port, set_signal_0_3_10_port, 
      set_signal_0_3_9_port, set_signal_0_3_8_port, set_signal_0_3_7_port, 
      set_signal_0_3_6_port, set_signal_0_3_5_port, set_signal_0_3_4_port, 
      set_signal_0_3_3_port, set_signal_0_3_2_port, set_signal_0_3_1_port, 
      set_signal_0_3_0_port, set_signal_0_4_15_port, set_signal_0_4_14_port, 
      set_signal_0_4_13_port, set_signal_0_4_12_port, set_signal_0_4_11_port, 
      set_signal_0_4_10_port, set_signal_0_4_9_port, set_signal_0_4_8_port, 
      set_signal_0_4_7_port, set_signal_0_4_6_port, set_signal_0_4_5_port, 
      set_signal_0_4_4_port, set_signal_0_4_3_port, set_signal_0_4_2_port, 
      set_signal_0_4_1_port, set_signal_0_4_0_port, set_signal_0_5_15_port, 
      set_signal_0_5_14_port, set_signal_0_5_13_port, set_signal_0_5_12_port, 
      set_signal_0_5_11_port, set_signal_0_5_10_port, set_signal_0_5_9_port, 
      set_signal_0_5_8_port, set_signal_0_5_7_port, set_signal_0_5_6_port, 
      set_signal_0_5_5_port, set_signal_0_5_4_port, set_signal_0_5_3_port, 
      set_signal_0_5_2_port, set_signal_0_5_1_port, set_signal_0_5_0_port, 
      set_signal_0_6_15_port, set_signal_0_6_14_port, set_signal_0_6_13_port, 
      set_signal_0_6_12_port, set_signal_0_6_11_port, set_signal_0_6_10_port, 
      set_signal_0_6_9_port, set_signal_0_6_8_port, set_signal_0_6_7_port, 
      set_signal_0_6_6_port, set_signal_0_6_5_port, set_signal_0_6_4_port, 
      set_signal_0_6_3_port, set_signal_0_6_2_port, set_signal_0_6_1_port, 
      set_signal_0_6_0_port, set_signal_1_1_15_port, set_signal_1_1_14_port, 
      set_signal_1_1_13_port, set_signal_1_1_12_port, set_signal_1_1_11_port, 
      set_signal_1_1_10_port, set_signal_1_1_9_port, set_signal_1_1_8_port, 
      set_signal_1_1_7_port, set_signal_1_1_6_port, set_signal_1_1_5_port, 
      set_signal_1_1_4_port, set_signal_1_1_3_port, set_signal_1_1_2_port, 
      set_signal_1_1_1_port, set_signal_1_1_0_port, set_signal_1_2_15_port, 
      set_signal_1_2_14_port, set_signal_1_2_13_port, set_signal_1_2_12_port, 
      set_signal_1_2_11_port, set_signal_1_2_10_port, set_signal_1_2_9_port, 
      set_signal_1_2_8_port, set_signal_1_2_7_port, set_signal_1_2_6_port, 
      set_signal_1_2_5_port, set_signal_1_2_4_port, set_signal_1_2_3_port, 
      set_signal_1_2_2_port, set_signal_1_2_1_port, set_signal_1_2_0_port, 
      set_signal_1_3_15_port, set_signal_1_3_14_port, set_signal_1_3_13_port, 
      set_signal_1_3_12_port, set_signal_1_3_11_port, set_signal_1_3_10_port, 
      set_signal_1_3_9_port, set_signal_1_3_8_port, set_signal_1_3_7_port, 
      set_signal_1_3_6_port, set_signal_1_3_5_port, set_signal_1_3_4_port, 
      set_signal_1_3_3_port, set_signal_1_3_2_port, set_signal_1_3_1_port, 
      set_signal_1_3_0_port, set_signal_1_4_15_port, set_signal_1_4_14_port, 
      set_signal_1_4_13_port, set_signal_1_4_12_port, set_signal_1_4_11_port, 
      set_signal_1_4_10_port, set_signal_1_4_9_port, set_signal_1_4_8_port, 
      set_signal_1_4_7_port, set_signal_1_4_6_port, set_signal_1_4_5_port, 
      set_signal_1_4_4_port, set_signal_1_4_3_port, set_signal_1_4_2_port, 
      set_signal_1_4_1_port, set_signal_1_4_0_port, set_signal_1_5_15_port, 
      set_signal_1_5_14_port, set_signal_1_5_13_port, set_signal_1_5_12_port, 
      set_signal_1_5_11_port, set_signal_1_5_10_port, set_signal_1_5_9_port, 
      set_signal_1_5_8_port, set_signal_1_5_7_port, set_signal_1_5_6_port, 
      set_signal_1_5_5_port, set_signal_1_5_4_port, set_signal_1_5_3_port, 
      set_signal_1_5_2_port, set_signal_1_5_1_port, set_signal_1_5_0_port, 
      set_signal_1_6_15_port, set_signal_1_6_14_port, set_signal_1_6_13_port, 
      set_signal_1_6_12_port, set_signal_1_6_11_port, set_signal_1_6_10_port, 
      set_signal_1_6_9_port, set_signal_1_6_8_port, set_signal_1_6_7_port, 
      set_signal_1_6_6_port, set_signal_1_6_5_port, set_signal_1_6_4_port, 
      set_signal_1_6_3_port, set_signal_1_6_2_port, set_signal_1_6_1_port, 
      set_signal_1_6_0_port, set_signal_2_1_15_port, set_signal_2_1_14_port, 
      set_signal_2_1_13_port, set_signal_2_1_12_port, set_signal_2_1_11_port, 
      set_signal_2_1_10_port, set_signal_2_1_9_port, set_signal_2_1_8_port, 
      set_signal_2_1_7_port, set_signal_2_1_6_port, set_signal_2_1_5_port, 
      set_signal_2_1_4_port, set_signal_2_1_3_port, set_signal_2_1_2_port, 
      set_signal_2_1_1_port, set_signal_2_1_0_port, set_signal_2_2_15_port, 
      set_signal_2_2_14_port, set_signal_2_2_13_port, set_signal_2_2_12_port, 
      set_signal_2_2_11_port, set_signal_2_2_10_port, set_signal_2_2_9_port, 
      set_signal_2_2_8_port, set_signal_2_2_7_port, set_signal_2_2_6_port, 
      set_signal_2_2_5_port, set_signal_2_2_4_port, set_signal_2_2_3_port, 
      set_signal_2_2_2_port, set_signal_2_2_1_port, set_signal_2_2_0_port, 
      set_signal_2_3_15_port, set_signal_2_3_14_port, set_signal_2_3_13_port, 
      set_signal_2_3_12_port, set_signal_2_3_11_port, set_signal_2_3_10_port, 
      set_signal_2_3_9_port, set_signal_2_3_8_port, set_signal_2_3_7_port, 
      set_signal_2_3_6_port, set_signal_2_3_5_port, set_signal_2_3_4_port, 
      set_signal_2_3_3_port, set_signal_2_3_2_port, set_signal_2_3_1_port, 
      set_signal_2_3_0_port, set_signal_2_4_15_port, set_signal_2_4_14_port, 
      set_signal_2_4_13_port, set_signal_2_4_12_port, set_signal_2_4_11_port, 
      set_signal_2_4_10_port, set_signal_2_4_9_port, set_signal_2_4_8_port, 
      set_signal_2_4_7_port, set_signal_2_4_6_port, set_signal_2_4_5_port, 
      set_signal_2_4_4_port, set_signal_2_4_3_port, set_signal_2_4_2_port, 
      set_signal_2_4_1_port, set_signal_2_4_0_port, set_signal_2_5_15_port, 
      set_signal_2_5_14_port, set_signal_2_5_13_port, set_signal_2_5_12_port, 
      set_signal_2_5_11_port, set_signal_2_5_10_port, set_signal_2_5_9_port, 
      set_signal_2_5_8_port, set_signal_2_5_7_port, set_signal_2_5_6_port, 
      set_signal_2_5_5_port, set_signal_2_5_4_port, set_signal_2_5_3_port, 
      set_signal_2_5_2_port, set_signal_2_5_1_port, set_signal_2_5_0_port, 
      set_signal_2_6_15_port, set_signal_2_6_14_port, set_signal_2_6_13_port, 
      set_signal_2_6_12_port, set_signal_2_6_11_port, set_signal_2_6_10_port, 
      set_signal_2_6_9_port, set_signal_2_6_8_port, set_signal_2_6_7_port, 
      set_signal_2_6_6_port, set_signal_2_6_5_port, set_signal_2_6_4_port, 
      set_signal_2_6_3_port, set_signal_2_6_2_port, set_signal_2_6_1_port, 
      set_signal_2_6_0_port, set_signal_3_1_15_port, set_signal_3_1_14_port, 
      set_signal_3_1_13_port, set_signal_3_1_12_port, set_signal_3_1_11_port, 
      set_signal_3_1_10_port, set_signal_3_1_9_port, set_signal_3_1_8_port, 
      set_signal_3_1_7_port, set_signal_3_1_6_port, set_signal_3_1_5_port, 
      set_signal_3_1_4_port, set_signal_3_1_3_port, set_signal_3_1_2_port, 
      set_signal_3_1_1_port, set_signal_3_1_0_port, set_signal_3_2_15_port, 
      set_signal_3_2_14_port, set_signal_3_2_13_port, set_signal_3_2_12_port, 
      set_signal_3_2_11_port, set_signal_3_2_10_port, set_signal_3_2_9_port, 
      set_signal_3_2_8_port, set_signal_3_2_7_port, set_signal_3_2_6_port, 
      set_signal_3_2_5_port, set_signal_3_2_4_port, set_signal_3_2_3_port, 
      set_signal_3_2_2_port, set_signal_3_2_1_port, set_signal_3_2_0_port, 
      set_signal_3_3_15_port, set_signal_3_3_14_port, set_signal_3_3_13_port, 
      set_signal_3_3_12_port, set_signal_3_3_11_port, set_signal_3_3_10_port, 
      set_signal_3_3_9_port, set_signal_3_3_8_port, set_signal_3_3_7_port, 
      set_signal_3_3_6_port, set_signal_3_3_5_port, set_signal_3_3_4_port, 
      set_signal_3_3_3_port, set_signal_3_3_2_port, set_signal_3_3_1_port, 
      set_signal_3_3_0_port, set_signal_3_4_15_port, set_signal_3_4_14_port, 
      set_signal_3_4_13_port, set_signal_3_4_12_port, set_signal_3_4_11_port, 
      set_signal_3_4_10_port, set_signal_3_4_9_port, set_signal_3_4_8_port, 
      set_signal_3_4_7_port, set_signal_3_4_6_port, set_signal_3_4_5_port, 
      set_signal_3_4_4_port, set_signal_3_4_3_port, set_signal_3_4_2_port, 
      set_signal_3_4_1_port, set_signal_3_4_0_port, set_signal_3_5_15_port, 
      set_signal_3_5_14_port, set_signal_3_5_13_port, set_signal_3_5_12_port, 
      set_signal_3_5_11_port, set_signal_3_5_10_port, set_signal_3_5_9_port, 
      set_signal_3_5_8_port, set_signal_3_5_7_port, set_signal_3_5_6_port, 
      set_signal_3_5_5_port, set_signal_3_5_4_port, set_signal_3_5_3_port, 
      set_signal_3_5_2_port, set_signal_3_5_1_port, set_signal_3_5_0_port, 
      enc_signal_0_1_2_port, enc_signal_0_1_1_port, enc_signal_0_1_0_port, 
      enc_signal_1_1_2_port, enc_signal_1_1_1_port, enc_signal_1_1_0_port, 
      enc_signal_2_1_2_port, enc_signal_2_1_1_port, enc_signal_2_1_0_port, 
      enc_signal_3_1_2_port, enc_signal_3_1_1_port, enc_signal_3_1_0_port, 
      rca_signal_1_0_15_port, rca_signal_1_0_14_port, rca_signal_1_0_13_port, 
      rca_signal_1_0_12_port, rca_signal_1_0_11_port, rca_signal_1_0_10_port, 
      rca_signal_1_0_9_port, rca_signal_1_0_8_port, rca_signal_1_0_7_port, 
      rca_signal_1_0_6_port, rca_signal_1_0_5_port, rca_signal_1_0_4_port, 
      rca_signal_1_0_3_port, rca_signal_1_0_2_port, rca_signal_1_0_1_port, 
      rca_signal_1_0_0_port, rca_signal_1_1_15_port, rca_signal_1_1_14_port, 
      rca_signal_1_1_13_port, rca_signal_1_1_12_port, rca_signal_1_1_11_port, 
      rca_signal_1_1_10_port, rca_signal_1_1_9_port, rca_signal_1_1_8_port, 
      rca_signal_1_1_7_port, rca_signal_1_1_6_port, rca_signal_1_1_5_port, 
      rca_signal_1_1_4_port, rca_signal_1_1_3_port, rca_signal_1_1_2_port, 
      rca_signal_1_1_1_port, rca_signal_1_1_0_port, rca_signal_2_0_15_port, 
      rca_signal_2_0_14_port, rca_signal_2_0_13_port, rca_signal_2_0_12_port, 
      rca_signal_2_0_11_port, rca_signal_2_0_10_port, rca_signal_2_0_9_port, 
      rca_signal_2_0_8_port, rca_signal_2_0_7_port, rca_signal_2_0_6_port, 
      rca_signal_2_0_5_port, rca_signal_2_0_4_port, rca_signal_2_0_3_port, 
      rca_signal_2_0_2_port, rca_signal_2_0_1_port, rca_signal_2_0_0_port, 
      rca_signal_2_1_15_port, rca_signal_2_1_14_port, rca_signal_2_1_13_port, 
      rca_signal_2_1_12_port, rca_signal_2_1_11_port, rca_signal_2_1_10_port, 
      rca_signal_2_1_9_port, rca_signal_2_1_8_port, rca_signal_2_1_7_port, 
      rca_signal_2_1_6_port, rca_signal_2_1_5_port, rca_signal_2_1_4_port, 
      rca_signal_2_1_3_port, rca_signal_2_1_2_port, rca_signal_2_1_1_port, 
      rca_signal_2_1_0_port, rca_signal_3_0_15_port, rca_signal_3_0_14_port, 
      rca_signal_3_0_13_port, rca_signal_3_0_12_port, rca_signal_3_0_11_port, 
      rca_signal_3_0_10_port, rca_signal_3_0_9_port, rca_signal_3_0_8_port, 
      rca_signal_3_0_7_port, rca_signal_3_0_6_port, rca_signal_3_0_5_port, 
      rca_signal_3_0_4_port, rca_signal_3_0_3_port, rca_signal_3_0_2_port, 
      rca_signal_3_0_1_port, rca_signal_3_0_0_port, rca_signal_3_1_15_port, 
      rca_signal_3_1_14_port, rca_signal_3_1_13_port, rca_signal_3_1_12_port, 
      rca_signal_3_1_11_port, rca_signal_3_1_10_port, rca_signal_3_1_9_port, 
      rca_signal_3_1_8_port, rca_signal_3_1_7_port, rca_signal_3_1_6_port, 
      rca_signal_3_1_5_port, rca_signal_3_1_4_port, rca_signal_3_1_3_port, 
      rca_signal_3_1_2_port, rca_signal_3_1_1_port, rca_signal_3_1_0_port, 
      n_1012, n_1013, n_1014, n_1015, n_1016, n_1017, n_1018, n_1019, n_1020, 
      n_1021, n_1022, n_1023, n_1024, n_1025, n_1026, n_1027, n_1028, n_1029, 
      n_1030, n_1031, n_1032, n_1033, n_1034, n_1035, n_1036, n_1037, n_1038, 
      n_1039, n_1040, n_1041, n_1042, n_1043, n_1044, n_1045, n_1046, n_1047, 
      n_1048, n_1049, n_1050, n_1051, n_1052, n_1053, n_1054, n_1055, n_1056, 
      n_1057, n_1058, n_1059, n_1060, n_1061, n_1062, n_1063, n_1064, n_1065, 
      n_1066, n_1067, n_1068, n_1069, n_1070, n_1071, n_1072, n_1073, n_1074, 
      n_1075, n_1076, n_1077, n_1078, n_1079, n_1080, n_1081, n_1082, n_1083, 
      n_1084, n_1085, n_1086, n_1087, n_1088, n_1089, n_1090, n_1091, n_1092, 
      n_1093, n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, n_1100, n_1101, 
      n_1102, n_1103, n_1104, n_1105, n_1106, n_1107, n_1108 : std_logic;

begin
   
   X_Logic0_port <= '0';
   enc0_0 : ENC3TO3_0 port map( X(2) => B_mp(1), X(1) => B_mp(0), X(0) => 
                           X_Logic0_port, Y(2) => enc_signal_0_1_2_port, Y(1) 
                           => enc_signal_0_1_1_port, Y(0) => 
                           enc_signal_0_1_0_port);
   set0_0 : SETTLER_NBIT16_0 port map( A(15) => A_mp(7), A(14) => A_mp(7), 
                           A(13) => A_mp(7), A(12) => A_mp(7), A(11) => A_mp(7)
                           , A(10) => A_mp(7), A(9) => A_mp(7), A(8) => A_mp(7)
                           , A(7) => A_mp(7), A(6) => A_mp(6), A(5) => A_mp(5),
                           A(4) => A_mp(4), A(3) => A_mp(3), A(2) => A_mp(2), 
                           A(1) => A_mp(1), A(0) => A_mp(0), Y0(15) => n_1012, 
                           Y0(14) => n_1013, Y0(13) => n_1014, Y0(12) => n_1015
                           , Y0(11) => n_1016, Y0(10) => n_1017, Y0(9) => 
                           n_1018, Y0(8) => n_1019, Y0(7) => n_1020, Y0(6) => 
                           n_1021, Y0(5) => n_1022, Y0(4) => n_1023, Y0(3) => 
                           n_1024, Y0(2) => n_1025, Y0(1) => n_1026, Y0(0) => 
                           n_1027, Y1(15) => set_signal_0_2_15_port, Y1(14) => 
                           set_signal_0_2_14_port, Y1(13) => 
                           set_signal_0_2_13_port, Y1(12) => 
                           set_signal_0_2_12_port, Y1(11) => 
                           set_signal_0_2_11_port, Y1(10) => 
                           set_signal_0_2_10_port, Y1(9) => 
                           set_signal_0_2_9_port, Y1(8) => 
                           set_signal_0_2_8_port, Y1(7) => 
                           set_signal_0_2_7_port, Y1(6) => 
                           set_signal_0_2_6_port, Y1(5) => 
                           set_signal_0_2_5_port, Y1(4) => 
                           set_signal_0_2_4_port, Y1(3) => 
                           set_signal_0_2_3_port, Y1(2) => 
                           set_signal_0_2_2_port, Y1(1) => 
                           set_signal_0_2_1_port, Y1(0) => 
                           set_signal_0_2_0_port, Y2(15) => 
                           set_signal_0_3_15_port, Y2(14) => 
                           set_signal_0_3_14_port, Y2(13) => 
                           set_signal_0_3_13_port, Y2(12) => 
                           set_signal_0_3_12_port, Y2(11) => 
                           set_signal_0_3_11_port, Y2(10) => 
                           set_signal_0_3_10_port, Y2(9) => 
                           set_signal_0_3_9_port, Y2(8) => 
                           set_signal_0_3_8_port, Y2(7) => 
                           set_signal_0_3_7_port, Y2(6) => 
                           set_signal_0_3_6_port, Y2(5) => 
                           set_signal_0_3_5_port, Y2(4) => 
                           set_signal_0_3_4_port, Y2(3) => 
                           set_signal_0_3_3_port, Y2(2) => 
                           set_signal_0_3_2_port, Y2(1) => 
                           set_signal_0_3_1_port, Y2(0) => 
                           set_signal_0_3_0_port, Y3(15) => 
                           set_signal_0_4_15_port, Y3(14) => 
                           set_signal_0_4_14_port, Y3(13) => 
                           set_signal_0_4_13_port, Y3(12) => 
                           set_signal_0_4_12_port, Y3(11) => 
                           set_signal_0_4_11_port, Y3(10) => 
                           set_signal_0_4_10_port, Y3(9) => 
                           set_signal_0_4_9_port, Y3(8) => 
                           set_signal_0_4_8_port, Y3(7) => 
                           set_signal_0_4_7_port, Y3(6) => 
                           set_signal_0_4_6_port, Y3(5) => 
                           set_signal_0_4_5_port, Y3(4) => 
                           set_signal_0_4_4_port, Y3(3) => 
                           set_signal_0_4_3_port, Y3(2) => 
                           set_signal_0_4_2_port, Y3(1) => 
                           set_signal_0_4_1_port, Y3(0) => n_1028, Y4(15) => 
                           set_signal_0_5_15_port, Y4(14) => 
                           set_signal_0_5_14_port, Y4(13) => 
                           set_signal_0_5_13_port, Y4(12) => 
                           set_signal_0_5_12_port, Y4(11) => 
                           set_signal_0_5_11_port, Y4(10) => 
                           set_signal_0_5_10_port, Y4(9) => 
                           set_signal_0_5_9_port, Y4(8) => 
                           set_signal_0_5_8_port, Y4(7) => 
                           set_signal_0_5_7_port, Y4(6) => 
                           set_signal_0_5_6_port, Y4(5) => 
                           set_signal_0_5_5_port, Y4(4) => 
                           set_signal_0_5_4_port, Y4(3) => 
                           set_signal_0_5_3_port, Y4(2) => 
                           set_signal_0_5_2_port, Y4(1) => 
                           set_signal_0_5_1_port, Y4(0) => n_1029, Y5(15) => 
                           set_signal_0_6_15_port, Y5(14) => 
                           set_signal_0_6_14_port, Y5(13) => 
                           set_signal_0_6_13_port, Y5(12) => 
                           set_signal_0_6_12_port, Y5(11) => 
                           set_signal_0_6_11_port, Y5(10) => 
                           set_signal_0_6_10_port, Y5(9) => 
                           set_signal_0_6_9_port, Y5(8) => 
                           set_signal_0_6_8_port, Y5(7) => 
                           set_signal_0_6_7_port, Y5(6) => 
                           set_signal_0_6_6_port, Y5(5) => 
                           set_signal_0_6_5_port, Y5(4) => 
                           set_signal_0_6_4_port, Y5(3) => 
                           set_signal_0_6_3_port, Y5(2) => 
                           set_signal_0_6_2_port, Y5(1) => n_1030, Y5(0) => 
                           n_1031);
   mux0_0 : MUX51_GENERIC_NBIT16_0 port map( A0(15) => set_signal_0_1_15_port, 
                           A0(14) => set_signal_0_1_14_port, A0(13) => 
                           set_signal_0_1_13_port, A0(12) => 
                           set_signal_0_1_12_port, A0(11) => 
                           set_signal_0_1_11_port, A0(10) => 
                           set_signal_0_1_10_port, A0(9) => 
                           set_signal_0_1_9_port, A0(8) => 
                           set_signal_0_1_8_port, A0(7) => 
                           set_signal_0_1_7_port, A0(6) => 
                           set_signal_0_1_6_port, A0(5) => 
                           set_signal_0_1_5_port, A0(4) => 
                           set_signal_0_1_4_port, A0(3) => 
                           set_signal_0_1_3_port, A0(2) => 
                           set_signal_0_1_2_port, A0(1) => 
                           set_signal_0_1_1_port, A0(0) => 
                           set_signal_0_1_0_port, A1(15) => 
                           set_signal_0_2_15_port, A1(14) => 
                           set_signal_0_2_14_port, A1(13) => 
                           set_signal_0_2_13_port, A1(12) => 
                           set_signal_0_2_12_port, A1(11) => 
                           set_signal_0_2_11_port, A1(10) => 
                           set_signal_0_2_10_port, A1(9) => 
                           set_signal_0_2_9_port, A1(8) => 
                           set_signal_0_2_8_port, A1(7) => 
                           set_signal_0_2_7_port, A1(6) => 
                           set_signal_0_2_6_port, A1(5) => 
                           set_signal_0_2_5_port, A1(4) => 
                           set_signal_0_2_4_port, A1(3) => 
                           set_signal_0_2_3_port, A1(2) => 
                           set_signal_0_2_2_port, A1(1) => 
                           set_signal_0_2_1_port, A1(0) => 
                           set_signal_0_2_0_port, A2(15) => 
                           set_signal_0_3_15_port, A2(14) => 
                           set_signal_0_3_14_port, A2(13) => 
                           set_signal_0_3_13_port, A2(12) => 
                           set_signal_0_3_12_port, A2(11) => 
                           set_signal_0_3_11_port, A2(10) => 
                           set_signal_0_3_10_port, A2(9) => 
                           set_signal_0_3_9_port, A2(8) => 
                           set_signal_0_3_8_port, A2(7) => 
                           set_signal_0_3_7_port, A2(6) => 
                           set_signal_0_3_6_port, A2(5) => 
                           set_signal_0_3_5_port, A2(4) => 
                           set_signal_0_3_4_port, A2(3) => 
                           set_signal_0_3_3_port, A2(2) => 
                           set_signal_0_3_2_port, A2(1) => 
                           set_signal_0_3_1_port, A2(0) => 
                           set_signal_0_3_0_port, A3(15) => 
                           set_signal_0_4_15_port, A3(14) => 
                           set_signal_0_4_14_port, A3(13) => 
                           set_signal_0_4_13_port, A3(12) => 
                           set_signal_0_4_12_port, A3(11) => 
                           set_signal_0_4_11_port, A3(10) => 
                           set_signal_0_4_10_port, A3(9) => 
                           set_signal_0_4_9_port, A3(8) => 
                           set_signal_0_4_8_port, A3(7) => 
                           set_signal_0_4_7_port, A3(6) => 
                           set_signal_0_4_6_port, A3(5) => 
                           set_signal_0_4_5_port, A3(4) => 
                           set_signal_0_4_4_port, A3(3) => 
                           set_signal_0_4_3_port, A3(2) => 
                           set_signal_0_4_2_port, A3(1) => 
                           set_signal_0_4_1_port, A3(0) => 
                           set_signal_0_4_0_port, A4(15) => 
                           set_signal_0_5_15_port, A4(14) => 
                           set_signal_0_5_14_port, A4(13) => 
                           set_signal_0_5_13_port, A4(12) => 
                           set_signal_0_5_12_port, A4(11) => 
                           set_signal_0_5_11_port, A4(10) => 
                           set_signal_0_5_10_port, A4(9) => 
                           set_signal_0_5_9_port, A4(8) => 
                           set_signal_0_5_8_port, A4(7) => 
                           set_signal_0_5_7_port, A4(6) => 
                           set_signal_0_5_6_port, A4(5) => 
                           set_signal_0_5_5_port, A4(4) => 
                           set_signal_0_5_4_port, A4(3) => 
                           set_signal_0_5_3_port, A4(2) => 
                           set_signal_0_5_2_port, A4(1) => 
                           set_signal_0_5_1_port, A4(0) => 
                           set_signal_0_5_0_port, SEL(2) => 
                           enc_signal_0_1_2_port, SEL(1) => 
                           enc_signal_0_1_1_port, SEL(0) => 
                           enc_signal_0_1_0_port, Y(15) => 
                           rca_signal_1_1_15_port, Y(14) => 
                           rca_signal_1_1_14_port, Y(13) => 
                           rca_signal_1_1_13_port, Y(12) => 
                           rca_signal_1_1_12_port, Y(11) => 
                           rca_signal_1_1_11_port, Y(10) => 
                           rca_signal_1_1_10_port, Y(9) => 
                           rca_signal_1_1_9_port, Y(8) => rca_signal_1_1_8_port
                           , Y(7) => rca_signal_1_1_7_port, Y(6) => 
                           rca_signal_1_1_6_port, Y(5) => rca_signal_1_1_5_port
                           , Y(4) => rca_signal_1_1_4_port, Y(3) => 
                           rca_signal_1_1_3_port, Y(2) => rca_signal_1_1_2_port
                           , Y(1) => rca_signal_1_1_1_port, Y(0) => 
                           rca_signal_1_1_0_port);
   enci_1 : ENC3TO3_3 port map( X(2) => B_mp(3), X(1) => B_mp(2), X(0) => 
                           B_mp(1), Y(2) => enc_signal_1_1_2_port, Y(1) => 
                           enc_signal_1_1_1_port, Y(0) => enc_signal_1_1_0_port
                           );
   seti_1 : SETTLER_NBIT16_3 port map( A(15) => set_signal_0_6_15_port, A(14) 
                           => set_signal_0_6_14_port, A(13) => 
                           set_signal_0_6_13_port, A(12) => 
                           set_signal_0_6_12_port, A(11) => 
                           set_signal_0_6_11_port, A(10) => 
                           set_signal_0_6_10_port, A(9) => 
                           set_signal_0_6_9_port, A(8) => set_signal_0_6_8_port
                           , A(7) => set_signal_0_6_7_port, A(6) => 
                           set_signal_0_6_6_port, A(5) => set_signal_0_6_5_port
                           , A(4) => set_signal_0_6_4_port, A(3) => 
                           set_signal_0_6_3_port, A(2) => set_signal_0_6_2_port
                           , A(1) => set_signal_0_6_1_port, A(0) => 
                           set_signal_0_6_0_port, Y0(15) => n_1032, Y0(14) => 
                           n_1033, Y0(13) => n_1034, Y0(12) => n_1035, Y0(11) 
                           => n_1036, Y0(10) => n_1037, Y0(9) => n_1038, Y0(8) 
                           => n_1039, Y0(7) => n_1040, Y0(6) => n_1041, Y0(5) 
                           => n_1042, Y0(4) => n_1043, Y0(3) => n_1044, Y0(2) 
                           => n_1045, Y0(1) => n_1046, Y0(0) => n_1047, Y1(15) 
                           => set_signal_1_2_15_port, Y1(14) => 
                           set_signal_1_2_14_port, Y1(13) => 
                           set_signal_1_2_13_port, Y1(12) => 
                           set_signal_1_2_12_port, Y1(11) => 
                           set_signal_1_2_11_port, Y1(10) => 
                           set_signal_1_2_10_port, Y1(9) => 
                           set_signal_1_2_9_port, Y1(8) => 
                           set_signal_1_2_8_port, Y1(7) => 
                           set_signal_1_2_7_port, Y1(6) => 
                           set_signal_1_2_6_port, Y1(5) => 
                           set_signal_1_2_5_port, Y1(4) => 
                           set_signal_1_2_4_port, Y1(3) => 
                           set_signal_1_2_3_port, Y1(2) => 
                           set_signal_1_2_2_port, Y1(1) => 
                           set_signal_1_2_1_port, Y1(0) => 
                           set_signal_1_2_0_port, Y2(15) => 
                           set_signal_1_3_15_port, Y2(14) => 
                           set_signal_1_3_14_port, Y2(13) => 
                           set_signal_1_3_13_port, Y2(12) => 
                           set_signal_1_3_12_port, Y2(11) => 
                           set_signal_1_3_11_port, Y2(10) => 
                           set_signal_1_3_10_port, Y2(9) => 
                           set_signal_1_3_9_port, Y2(8) => 
                           set_signal_1_3_8_port, Y2(7) => 
                           set_signal_1_3_7_port, Y2(6) => 
                           set_signal_1_3_6_port, Y2(5) => 
                           set_signal_1_3_5_port, Y2(4) => 
                           set_signal_1_3_4_port, Y2(3) => 
                           set_signal_1_3_3_port, Y2(2) => 
                           set_signal_1_3_2_port, Y2(1) => 
                           set_signal_1_3_1_port, Y2(0) => 
                           set_signal_1_3_0_port, Y3(15) => 
                           set_signal_1_4_15_port, Y3(14) => 
                           set_signal_1_4_14_port, Y3(13) => 
                           set_signal_1_4_13_port, Y3(12) => 
                           set_signal_1_4_12_port, Y3(11) => 
                           set_signal_1_4_11_port, Y3(10) => 
                           set_signal_1_4_10_port, Y3(9) => 
                           set_signal_1_4_9_port, Y3(8) => 
                           set_signal_1_4_8_port, Y3(7) => 
                           set_signal_1_4_7_port, Y3(6) => 
                           set_signal_1_4_6_port, Y3(5) => 
                           set_signal_1_4_5_port, Y3(4) => 
                           set_signal_1_4_4_port, Y3(3) => 
                           set_signal_1_4_3_port, Y3(2) => 
                           set_signal_1_4_2_port, Y3(1) => 
                           set_signal_1_4_1_port, Y3(0) => n_1048, Y4(15) => 
                           set_signal_1_5_15_port, Y4(14) => 
                           set_signal_1_5_14_port, Y4(13) => 
                           set_signal_1_5_13_port, Y4(12) => 
                           set_signal_1_5_12_port, Y4(11) => 
                           set_signal_1_5_11_port, Y4(10) => 
                           set_signal_1_5_10_port, Y4(9) => 
                           set_signal_1_5_9_port, Y4(8) => 
                           set_signal_1_5_8_port, Y4(7) => 
                           set_signal_1_5_7_port, Y4(6) => 
                           set_signal_1_5_6_port, Y4(5) => 
                           set_signal_1_5_5_port, Y4(4) => 
                           set_signal_1_5_4_port, Y4(3) => 
                           set_signal_1_5_3_port, Y4(2) => 
                           set_signal_1_5_2_port, Y4(1) => 
                           set_signal_1_5_1_port, Y4(0) => n_1049, Y5(15) => 
                           set_signal_1_6_15_port, Y5(14) => 
                           set_signal_1_6_14_port, Y5(13) => 
                           set_signal_1_6_13_port, Y5(12) => 
                           set_signal_1_6_12_port, Y5(11) => 
                           set_signal_1_6_11_port, Y5(10) => 
                           set_signal_1_6_10_port, Y5(9) => 
                           set_signal_1_6_9_port, Y5(8) => 
                           set_signal_1_6_8_port, Y5(7) => 
                           set_signal_1_6_7_port, Y5(6) => 
                           set_signal_1_6_6_port, Y5(5) => 
                           set_signal_1_6_5_port, Y5(4) => 
                           set_signal_1_6_4_port, Y5(3) => 
                           set_signal_1_6_3_port, Y5(2) => 
                           set_signal_1_6_2_port, Y5(1) => n_1050, Y5(0) => 
                           n_1051);
   muxi_1 : MUX51_GENERIC_NBIT16_3 port map( A0(15) => set_signal_1_1_15_port, 
                           A0(14) => set_signal_1_1_14_port, A0(13) => 
                           set_signal_1_1_13_port, A0(12) => 
                           set_signal_1_1_12_port, A0(11) => 
                           set_signal_1_1_11_port, A0(10) => 
                           set_signal_1_1_10_port, A0(9) => 
                           set_signal_1_1_9_port, A0(8) => 
                           set_signal_1_1_8_port, A0(7) => 
                           set_signal_1_1_7_port, A0(6) => 
                           set_signal_1_1_6_port, A0(5) => 
                           set_signal_1_1_5_port, A0(4) => 
                           set_signal_1_1_4_port, A0(3) => 
                           set_signal_1_1_3_port, A0(2) => 
                           set_signal_1_1_2_port, A0(1) => 
                           set_signal_1_1_1_port, A0(0) => 
                           set_signal_1_1_0_port, A1(15) => 
                           set_signal_1_2_15_port, A1(14) => 
                           set_signal_1_2_14_port, A1(13) => 
                           set_signal_1_2_13_port, A1(12) => 
                           set_signal_1_2_12_port, A1(11) => 
                           set_signal_1_2_11_port, A1(10) => 
                           set_signal_1_2_10_port, A1(9) => 
                           set_signal_1_2_9_port, A1(8) => 
                           set_signal_1_2_8_port, A1(7) => 
                           set_signal_1_2_7_port, A1(6) => 
                           set_signal_1_2_6_port, A1(5) => 
                           set_signal_1_2_5_port, A1(4) => 
                           set_signal_1_2_4_port, A1(3) => 
                           set_signal_1_2_3_port, A1(2) => 
                           set_signal_1_2_2_port, A1(1) => 
                           set_signal_1_2_1_port, A1(0) => 
                           set_signal_1_2_0_port, A2(15) => 
                           set_signal_1_3_15_port, A2(14) => 
                           set_signal_1_3_14_port, A2(13) => 
                           set_signal_1_3_13_port, A2(12) => 
                           set_signal_1_3_12_port, A2(11) => 
                           set_signal_1_3_11_port, A2(10) => 
                           set_signal_1_3_10_port, A2(9) => 
                           set_signal_1_3_9_port, A2(8) => 
                           set_signal_1_3_8_port, A2(7) => 
                           set_signal_1_3_7_port, A2(6) => 
                           set_signal_1_3_6_port, A2(5) => 
                           set_signal_1_3_5_port, A2(4) => 
                           set_signal_1_3_4_port, A2(3) => 
                           set_signal_1_3_3_port, A2(2) => 
                           set_signal_1_3_2_port, A2(1) => 
                           set_signal_1_3_1_port, A2(0) => 
                           set_signal_1_3_0_port, A3(15) => 
                           set_signal_1_4_15_port, A3(14) => 
                           set_signal_1_4_14_port, A3(13) => 
                           set_signal_1_4_13_port, A3(12) => 
                           set_signal_1_4_12_port, A3(11) => 
                           set_signal_1_4_11_port, A3(10) => 
                           set_signal_1_4_10_port, A3(9) => 
                           set_signal_1_4_9_port, A3(8) => 
                           set_signal_1_4_8_port, A3(7) => 
                           set_signal_1_4_7_port, A3(6) => 
                           set_signal_1_4_6_port, A3(5) => 
                           set_signal_1_4_5_port, A3(4) => 
                           set_signal_1_4_4_port, A3(3) => 
                           set_signal_1_4_3_port, A3(2) => 
                           set_signal_1_4_2_port, A3(1) => 
                           set_signal_1_4_1_port, A3(0) => 
                           set_signal_1_4_0_port, A4(15) => 
                           set_signal_1_5_15_port, A4(14) => 
                           set_signal_1_5_14_port, A4(13) => 
                           set_signal_1_5_13_port, A4(12) => 
                           set_signal_1_5_12_port, A4(11) => 
                           set_signal_1_5_11_port, A4(10) => 
                           set_signal_1_5_10_port, A4(9) => 
                           set_signal_1_5_9_port, A4(8) => 
                           set_signal_1_5_8_port, A4(7) => 
                           set_signal_1_5_7_port, A4(6) => 
                           set_signal_1_5_6_port, A4(5) => 
                           set_signal_1_5_5_port, A4(4) => 
                           set_signal_1_5_4_port, A4(3) => 
                           set_signal_1_5_3_port, A4(2) => 
                           set_signal_1_5_2_port, A4(1) => 
                           set_signal_1_5_1_port, A4(0) => 
                           set_signal_1_5_0_port, SEL(2) => 
                           enc_signal_1_1_2_port, SEL(1) => 
                           enc_signal_1_1_1_port, SEL(0) => 
                           enc_signal_1_1_0_port, Y(15) => 
                           rca_signal_1_0_15_port, Y(14) => 
                           rca_signal_1_0_14_port, Y(13) => 
                           rca_signal_1_0_13_port, Y(12) => 
                           rca_signal_1_0_12_port, Y(11) => 
                           rca_signal_1_0_11_port, Y(10) => 
                           rca_signal_1_0_10_port, Y(9) => 
                           rca_signal_1_0_9_port, Y(8) => rca_signal_1_0_8_port
                           , Y(7) => rca_signal_1_0_7_port, Y(6) => 
                           rca_signal_1_0_6_port, Y(5) => rca_signal_1_0_5_port
                           , Y(4) => rca_signal_1_0_4_port, Y(3) => 
                           rca_signal_1_0_3_port, Y(2) => rca_signal_1_0_2_port
                           , Y(1) => rca_signal_1_0_1_port, Y(0) => 
                           rca_signal_1_0_0_port);
   rcai_1 : RCA_size16_0 port map( a(15) => rca_signal_1_0_15_port, a(14) => 
                           rca_signal_1_0_14_port, a(13) => 
                           rca_signal_1_0_13_port, a(12) => 
                           rca_signal_1_0_12_port, a(11) => 
                           rca_signal_1_0_11_port, a(10) => 
                           rca_signal_1_0_10_port, a(9) => 
                           rca_signal_1_0_9_port, a(8) => rca_signal_1_0_8_port
                           , a(7) => rca_signal_1_0_7_port, a(6) => 
                           rca_signal_1_0_6_port, a(5) => rca_signal_1_0_5_port
                           , a(4) => rca_signal_1_0_4_port, a(3) => 
                           rca_signal_1_0_3_port, a(2) => rca_signal_1_0_2_port
                           , a(1) => rca_signal_1_0_1_port, a(0) => 
                           rca_signal_1_0_0_port, b(15) => 
                           rca_signal_1_1_15_port, b(14) => 
                           rca_signal_1_1_14_port, b(13) => 
                           rca_signal_1_1_13_port, b(12) => 
                           rca_signal_1_1_12_port, b(11) => 
                           rca_signal_1_1_11_port, b(10) => 
                           rca_signal_1_1_10_port, b(9) => 
                           rca_signal_1_1_9_port, b(8) => rca_signal_1_1_8_port
                           , b(7) => rca_signal_1_1_7_port, b(6) => 
                           rca_signal_1_1_6_port, b(5) => rca_signal_1_1_5_port
                           , b(4) => rca_signal_1_1_4_port, b(3) => 
                           rca_signal_1_1_3_port, b(2) => rca_signal_1_1_2_port
                           , b(1) => rca_signal_1_1_1_port, b(0) => 
                           rca_signal_1_1_0_port, c_in => X_Logic0_port, c_out 
                           => n_1052, sum(15) => rca_signal_2_1_15_port, 
                           sum(14) => rca_signal_2_1_14_port, sum(13) => 
                           rca_signal_2_1_13_port, sum(12) => 
                           rca_signal_2_1_12_port, sum(11) => 
                           rca_signal_2_1_11_port, sum(10) => 
                           rca_signal_2_1_10_port, sum(9) => 
                           rca_signal_2_1_9_port, sum(8) => 
                           rca_signal_2_1_8_port, sum(7) => 
                           rca_signal_2_1_7_port, sum(6) => 
                           rca_signal_2_1_6_port, sum(5) => 
                           rca_signal_2_1_5_port, sum(4) => 
                           rca_signal_2_1_4_port, sum(3) => 
                           rca_signal_2_1_3_port, sum(2) => 
                           rca_signal_2_1_2_port, sum(1) => 
                           rca_signal_2_1_1_port, sum(0) => 
                           rca_signal_2_1_0_port);
   enci_2 : ENC3TO3_2 port map( X(2) => B_mp(5), X(1) => B_mp(4), X(0) => 
                           B_mp(3), Y(2) => enc_signal_2_1_2_port, Y(1) => 
                           enc_signal_2_1_1_port, Y(0) => enc_signal_2_1_0_port
                           );
   seti_2 : SETTLER_NBIT16_2 port map( A(15) => set_signal_1_6_15_port, A(14) 
                           => set_signal_1_6_14_port, A(13) => 
                           set_signal_1_6_13_port, A(12) => 
                           set_signal_1_6_12_port, A(11) => 
                           set_signal_1_6_11_port, A(10) => 
                           set_signal_1_6_10_port, A(9) => 
                           set_signal_1_6_9_port, A(8) => set_signal_1_6_8_port
                           , A(7) => set_signal_1_6_7_port, A(6) => 
                           set_signal_1_6_6_port, A(5) => set_signal_1_6_5_port
                           , A(4) => set_signal_1_6_4_port, A(3) => 
                           set_signal_1_6_3_port, A(2) => set_signal_1_6_2_port
                           , A(1) => set_signal_1_6_1_port, A(0) => 
                           set_signal_1_6_0_port, Y0(15) => n_1053, Y0(14) => 
                           n_1054, Y0(13) => n_1055, Y0(12) => n_1056, Y0(11) 
                           => n_1057, Y0(10) => n_1058, Y0(9) => n_1059, Y0(8) 
                           => n_1060, Y0(7) => n_1061, Y0(6) => n_1062, Y0(5) 
                           => n_1063, Y0(4) => n_1064, Y0(3) => n_1065, Y0(2) 
                           => n_1066, Y0(1) => n_1067, Y0(0) => n_1068, Y1(15) 
                           => set_signal_2_2_15_port, Y1(14) => 
                           set_signal_2_2_14_port, Y1(13) => 
                           set_signal_2_2_13_port, Y1(12) => 
                           set_signal_2_2_12_port, Y1(11) => 
                           set_signal_2_2_11_port, Y1(10) => 
                           set_signal_2_2_10_port, Y1(9) => 
                           set_signal_2_2_9_port, Y1(8) => 
                           set_signal_2_2_8_port, Y1(7) => 
                           set_signal_2_2_7_port, Y1(6) => 
                           set_signal_2_2_6_port, Y1(5) => 
                           set_signal_2_2_5_port, Y1(4) => 
                           set_signal_2_2_4_port, Y1(3) => 
                           set_signal_2_2_3_port, Y1(2) => 
                           set_signal_2_2_2_port, Y1(1) => 
                           set_signal_2_2_1_port, Y1(0) => 
                           set_signal_2_2_0_port, Y2(15) => 
                           set_signal_2_3_15_port, Y2(14) => 
                           set_signal_2_3_14_port, Y2(13) => 
                           set_signal_2_3_13_port, Y2(12) => 
                           set_signal_2_3_12_port, Y2(11) => 
                           set_signal_2_3_11_port, Y2(10) => 
                           set_signal_2_3_10_port, Y2(9) => 
                           set_signal_2_3_9_port, Y2(8) => 
                           set_signal_2_3_8_port, Y2(7) => 
                           set_signal_2_3_7_port, Y2(6) => 
                           set_signal_2_3_6_port, Y2(5) => 
                           set_signal_2_3_5_port, Y2(4) => 
                           set_signal_2_3_4_port, Y2(3) => 
                           set_signal_2_3_3_port, Y2(2) => 
                           set_signal_2_3_2_port, Y2(1) => 
                           set_signal_2_3_1_port, Y2(0) => 
                           set_signal_2_3_0_port, Y3(15) => 
                           set_signal_2_4_15_port, Y3(14) => 
                           set_signal_2_4_14_port, Y3(13) => 
                           set_signal_2_4_13_port, Y3(12) => 
                           set_signal_2_4_12_port, Y3(11) => 
                           set_signal_2_4_11_port, Y3(10) => 
                           set_signal_2_4_10_port, Y3(9) => 
                           set_signal_2_4_9_port, Y3(8) => 
                           set_signal_2_4_8_port, Y3(7) => 
                           set_signal_2_4_7_port, Y3(6) => 
                           set_signal_2_4_6_port, Y3(5) => 
                           set_signal_2_4_5_port, Y3(4) => 
                           set_signal_2_4_4_port, Y3(3) => 
                           set_signal_2_4_3_port, Y3(2) => 
                           set_signal_2_4_2_port, Y3(1) => 
                           set_signal_2_4_1_port, Y3(0) => n_1069, Y4(15) => 
                           set_signal_2_5_15_port, Y4(14) => 
                           set_signal_2_5_14_port, Y4(13) => 
                           set_signal_2_5_13_port, Y4(12) => 
                           set_signal_2_5_12_port, Y4(11) => 
                           set_signal_2_5_11_port, Y4(10) => 
                           set_signal_2_5_10_port, Y4(9) => 
                           set_signal_2_5_9_port, Y4(8) => 
                           set_signal_2_5_8_port, Y4(7) => 
                           set_signal_2_5_7_port, Y4(6) => 
                           set_signal_2_5_6_port, Y4(5) => 
                           set_signal_2_5_5_port, Y4(4) => 
                           set_signal_2_5_4_port, Y4(3) => 
                           set_signal_2_5_3_port, Y4(2) => 
                           set_signal_2_5_2_port, Y4(1) => 
                           set_signal_2_5_1_port, Y4(0) => n_1070, Y5(15) => 
                           set_signal_2_6_15_port, Y5(14) => 
                           set_signal_2_6_14_port, Y5(13) => 
                           set_signal_2_6_13_port, Y5(12) => 
                           set_signal_2_6_12_port, Y5(11) => 
                           set_signal_2_6_11_port, Y5(10) => 
                           set_signal_2_6_10_port, Y5(9) => 
                           set_signal_2_6_9_port, Y5(8) => 
                           set_signal_2_6_8_port, Y5(7) => 
                           set_signal_2_6_7_port, Y5(6) => 
                           set_signal_2_6_6_port, Y5(5) => 
                           set_signal_2_6_5_port, Y5(4) => 
                           set_signal_2_6_4_port, Y5(3) => 
                           set_signal_2_6_3_port, Y5(2) => 
                           set_signal_2_6_2_port, Y5(1) => n_1071, Y5(0) => 
                           n_1072);
   muxi_2 : MUX51_GENERIC_NBIT16_2 port map( A0(15) => set_signal_2_1_15_port, 
                           A0(14) => set_signal_2_1_14_port, A0(13) => 
                           set_signal_2_1_13_port, A0(12) => 
                           set_signal_2_1_12_port, A0(11) => 
                           set_signal_2_1_11_port, A0(10) => 
                           set_signal_2_1_10_port, A0(9) => 
                           set_signal_2_1_9_port, A0(8) => 
                           set_signal_2_1_8_port, A0(7) => 
                           set_signal_2_1_7_port, A0(6) => 
                           set_signal_2_1_6_port, A0(5) => 
                           set_signal_2_1_5_port, A0(4) => 
                           set_signal_2_1_4_port, A0(3) => 
                           set_signal_2_1_3_port, A0(2) => 
                           set_signal_2_1_2_port, A0(1) => 
                           set_signal_2_1_1_port, A0(0) => 
                           set_signal_2_1_0_port, A1(15) => 
                           set_signal_2_2_15_port, A1(14) => 
                           set_signal_2_2_14_port, A1(13) => 
                           set_signal_2_2_13_port, A1(12) => 
                           set_signal_2_2_12_port, A1(11) => 
                           set_signal_2_2_11_port, A1(10) => 
                           set_signal_2_2_10_port, A1(9) => 
                           set_signal_2_2_9_port, A1(8) => 
                           set_signal_2_2_8_port, A1(7) => 
                           set_signal_2_2_7_port, A1(6) => 
                           set_signal_2_2_6_port, A1(5) => 
                           set_signal_2_2_5_port, A1(4) => 
                           set_signal_2_2_4_port, A1(3) => 
                           set_signal_2_2_3_port, A1(2) => 
                           set_signal_2_2_2_port, A1(1) => 
                           set_signal_2_2_1_port, A1(0) => 
                           set_signal_2_2_0_port, A2(15) => 
                           set_signal_2_3_15_port, A2(14) => 
                           set_signal_2_3_14_port, A2(13) => 
                           set_signal_2_3_13_port, A2(12) => 
                           set_signal_2_3_12_port, A2(11) => 
                           set_signal_2_3_11_port, A2(10) => 
                           set_signal_2_3_10_port, A2(9) => 
                           set_signal_2_3_9_port, A2(8) => 
                           set_signal_2_3_8_port, A2(7) => 
                           set_signal_2_3_7_port, A2(6) => 
                           set_signal_2_3_6_port, A2(5) => 
                           set_signal_2_3_5_port, A2(4) => 
                           set_signal_2_3_4_port, A2(3) => 
                           set_signal_2_3_3_port, A2(2) => 
                           set_signal_2_3_2_port, A2(1) => 
                           set_signal_2_3_1_port, A2(0) => 
                           set_signal_2_3_0_port, A3(15) => 
                           set_signal_2_4_15_port, A3(14) => 
                           set_signal_2_4_14_port, A3(13) => 
                           set_signal_2_4_13_port, A3(12) => 
                           set_signal_2_4_12_port, A3(11) => 
                           set_signal_2_4_11_port, A3(10) => 
                           set_signal_2_4_10_port, A3(9) => 
                           set_signal_2_4_9_port, A3(8) => 
                           set_signal_2_4_8_port, A3(7) => 
                           set_signal_2_4_7_port, A3(6) => 
                           set_signal_2_4_6_port, A3(5) => 
                           set_signal_2_4_5_port, A3(4) => 
                           set_signal_2_4_4_port, A3(3) => 
                           set_signal_2_4_3_port, A3(2) => 
                           set_signal_2_4_2_port, A3(1) => 
                           set_signal_2_4_1_port, A3(0) => 
                           set_signal_2_4_0_port, A4(15) => 
                           set_signal_2_5_15_port, A4(14) => 
                           set_signal_2_5_14_port, A4(13) => 
                           set_signal_2_5_13_port, A4(12) => 
                           set_signal_2_5_12_port, A4(11) => 
                           set_signal_2_5_11_port, A4(10) => 
                           set_signal_2_5_10_port, A4(9) => 
                           set_signal_2_5_9_port, A4(8) => 
                           set_signal_2_5_8_port, A4(7) => 
                           set_signal_2_5_7_port, A4(6) => 
                           set_signal_2_5_6_port, A4(5) => 
                           set_signal_2_5_5_port, A4(4) => 
                           set_signal_2_5_4_port, A4(3) => 
                           set_signal_2_5_3_port, A4(2) => 
                           set_signal_2_5_2_port, A4(1) => 
                           set_signal_2_5_1_port, A4(0) => 
                           set_signal_2_5_0_port, SEL(2) => 
                           enc_signal_2_1_2_port, SEL(1) => 
                           enc_signal_2_1_1_port, SEL(0) => 
                           enc_signal_2_1_0_port, Y(15) => 
                           rca_signal_2_0_15_port, Y(14) => 
                           rca_signal_2_0_14_port, Y(13) => 
                           rca_signal_2_0_13_port, Y(12) => 
                           rca_signal_2_0_12_port, Y(11) => 
                           rca_signal_2_0_11_port, Y(10) => 
                           rca_signal_2_0_10_port, Y(9) => 
                           rca_signal_2_0_9_port, Y(8) => rca_signal_2_0_8_port
                           , Y(7) => rca_signal_2_0_7_port, Y(6) => 
                           rca_signal_2_0_6_port, Y(5) => rca_signal_2_0_5_port
                           , Y(4) => rca_signal_2_0_4_port, Y(3) => 
                           rca_signal_2_0_3_port, Y(2) => rca_signal_2_0_2_port
                           , Y(1) => rca_signal_2_0_1_port, Y(0) => 
                           rca_signal_2_0_0_port);
   rcai_2 : RCA_size16_2 port map( a(15) => rca_signal_2_0_15_port, a(14) => 
                           rca_signal_2_0_14_port, a(13) => 
                           rca_signal_2_0_13_port, a(12) => 
                           rca_signal_2_0_12_port, a(11) => 
                           rca_signal_2_0_11_port, a(10) => 
                           rca_signal_2_0_10_port, a(9) => 
                           rca_signal_2_0_9_port, a(8) => rca_signal_2_0_8_port
                           , a(7) => rca_signal_2_0_7_port, a(6) => 
                           rca_signal_2_0_6_port, a(5) => rca_signal_2_0_5_port
                           , a(4) => rca_signal_2_0_4_port, a(3) => 
                           rca_signal_2_0_3_port, a(2) => rca_signal_2_0_2_port
                           , a(1) => rca_signal_2_0_1_port, a(0) => 
                           rca_signal_2_0_0_port, b(15) => 
                           rca_signal_2_1_15_port, b(14) => 
                           rca_signal_2_1_14_port, b(13) => 
                           rca_signal_2_1_13_port, b(12) => 
                           rca_signal_2_1_12_port, b(11) => 
                           rca_signal_2_1_11_port, b(10) => 
                           rca_signal_2_1_10_port, b(9) => 
                           rca_signal_2_1_9_port, b(8) => rca_signal_2_1_8_port
                           , b(7) => rca_signal_2_1_7_port, b(6) => 
                           rca_signal_2_1_6_port, b(5) => rca_signal_2_1_5_port
                           , b(4) => rca_signal_2_1_4_port, b(3) => 
                           rca_signal_2_1_3_port, b(2) => rca_signal_2_1_2_port
                           , b(1) => rca_signal_2_1_1_port, b(0) => 
                           rca_signal_2_1_0_port, c_in => X_Logic0_port, c_out 
                           => n_1073, sum(15) => rca_signal_3_1_15_port, 
                           sum(14) => rca_signal_3_1_14_port, sum(13) => 
                           rca_signal_3_1_13_port, sum(12) => 
                           rca_signal_3_1_12_port, sum(11) => 
                           rca_signal_3_1_11_port, sum(10) => 
                           rca_signal_3_1_10_port, sum(9) => 
                           rca_signal_3_1_9_port, sum(8) => 
                           rca_signal_3_1_8_port, sum(7) => 
                           rca_signal_3_1_7_port, sum(6) => 
                           rca_signal_3_1_6_port, sum(5) => 
                           rca_signal_3_1_5_port, sum(4) => 
                           rca_signal_3_1_4_port, sum(3) => 
                           rca_signal_3_1_3_port, sum(2) => 
                           rca_signal_3_1_2_port, sum(1) => 
                           rca_signal_3_1_1_port, sum(0) => 
                           rca_signal_3_1_0_port);
   enci_3 : ENC3TO3_1 port map( X(2) => B_mp(7), X(1) => B_mp(6), X(0) => 
                           B_mp(5), Y(2) => enc_signal_3_1_2_port, Y(1) => 
                           enc_signal_3_1_1_port, Y(0) => enc_signal_3_1_0_port
                           );
   seti_3 : SETTLER_NBIT16_1 port map( A(15) => set_signal_2_6_15_port, A(14) 
                           => set_signal_2_6_14_port, A(13) => 
                           set_signal_2_6_13_port, A(12) => 
                           set_signal_2_6_12_port, A(11) => 
                           set_signal_2_6_11_port, A(10) => 
                           set_signal_2_6_10_port, A(9) => 
                           set_signal_2_6_9_port, A(8) => set_signal_2_6_8_port
                           , A(7) => set_signal_2_6_7_port, A(6) => 
                           set_signal_2_6_6_port, A(5) => set_signal_2_6_5_port
                           , A(4) => set_signal_2_6_4_port, A(3) => 
                           set_signal_2_6_3_port, A(2) => set_signal_2_6_2_port
                           , A(1) => set_signal_2_6_1_port, A(0) => 
                           set_signal_2_6_0_port, Y0(15) => n_1074, Y0(14) => 
                           n_1075, Y0(13) => n_1076, Y0(12) => n_1077, Y0(11) 
                           => n_1078, Y0(10) => n_1079, Y0(9) => n_1080, Y0(8) 
                           => n_1081, Y0(7) => n_1082, Y0(6) => n_1083, Y0(5) 
                           => n_1084, Y0(4) => n_1085, Y0(3) => n_1086, Y0(2) 
                           => n_1087, Y0(1) => n_1088, Y0(0) => n_1089, Y1(15) 
                           => set_signal_3_2_15_port, Y1(14) => 
                           set_signal_3_2_14_port, Y1(13) => 
                           set_signal_3_2_13_port, Y1(12) => 
                           set_signal_3_2_12_port, Y1(11) => 
                           set_signal_3_2_11_port, Y1(10) => 
                           set_signal_3_2_10_port, Y1(9) => 
                           set_signal_3_2_9_port, Y1(8) => 
                           set_signal_3_2_8_port, Y1(7) => 
                           set_signal_3_2_7_port, Y1(6) => 
                           set_signal_3_2_6_port, Y1(5) => 
                           set_signal_3_2_5_port, Y1(4) => 
                           set_signal_3_2_4_port, Y1(3) => 
                           set_signal_3_2_3_port, Y1(2) => 
                           set_signal_3_2_2_port, Y1(1) => 
                           set_signal_3_2_1_port, Y1(0) => 
                           set_signal_3_2_0_port, Y2(15) => 
                           set_signal_3_3_15_port, Y2(14) => 
                           set_signal_3_3_14_port, Y2(13) => 
                           set_signal_3_3_13_port, Y2(12) => 
                           set_signal_3_3_12_port, Y2(11) => 
                           set_signal_3_3_11_port, Y2(10) => 
                           set_signal_3_3_10_port, Y2(9) => 
                           set_signal_3_3_9_port, Y2(8) => 
                           set_signal_3_3_8_port, Y2(7) => 
                           set_signal_3_3_7_port, Y2(6) => 
                           set_signal_3_3_6_port, Y2(5) => 
                           set_signal_3_3_5_port, Y2(4) => 
                           set_signal_3_3_4_port, Y2(3) => 
                           set_signal_3_3_3_port, Y2(2) => 
                           set_signal_3_3_2_port, Y2(1) => 
                           set_signal_3_3_1_port, Y2(0) => 
                           set_signal_3_3_0_port, Y3(15) => 
                           set_signal_3_4_15_port, Y3(14) => 
                           set_signal_3_4_14_port, Y3(13) => 
                           set_signal_3_4_13_port, Y3(12) => 
                           set_signal_3_4_12_port, Y3(11) => 
                           set_signal_3_4_11_port, Y3(10) => 
                           set_signal_3_4_10_port, Y3(9) => 
                           set_signal_3_4_9_port, Y3(8) => 
                           set_signal_3_4_8_port, Y3(7) => 
                           set_signal_3_4_7_port, Y3(6) => 
                           set_signal_3_4_6_port, Y3(5) => 
                           set_signal_3_4_5_port, Y3(4) => 
                           set_signal_3_4_4_port, Y3(3) => 
                           set_signal_3_4_3_port, Y3(2) => 
                           set_signal_3_4_2_port, Y3(1) => 
                           set_signal_3_4_1_port, Y3(0) => n_1090, Y4(15) => 
                           set_signal_3_5_15_port, Y4(14) => 
                           set_signal_3_5_14_port, Y4(13) => 
                           set_signal_3_5_13_port, Y4(12) => 
                           set_signal_3_5_12_port, Y4(11) => 
                           set_signal_3_5_11_port, Y4(10) => 
                           set_signal_3_5_10_port, Y4(9) => 
                           set_signal_3_5_9_port, Y4(8) => 
                           set_signal_3_5_8_port, Y4(7) => 
                           set_signal_3_5_7_port, Y4(6) => 
                           set_signal_3_5_6_port, Y4(5) => 
                           set_signal_3_5_5_port, Y4(4) => 
                           set_signal_3_5_4_port, Y4(3) => 
                           set_signal_3_5_3_port, Y4(2) => 
                           set_signal_3_5_2_port, Y4(1) => 
                           set_signal_3_5_1_port, Y4(0) => n_1091, Y5(15) => 
                           n_1092, Y5(14) => n_1093, Y5(13) => n_1094, Y5(12) 
                           => n_1095, Y5(11) => n_1096, Y5(10) => n_1097, Y5(9)
                           => n_1098, Y5(8) => n_1099, Y5(7) => n_1100, Y5(6) 
                           => n_1101, Y5(5) => n_1102, Y5(4) => n_1103, Y5(3) 
                           => n_1104, Y5(2) => n_1105, Y5(1) => n_1106, Y5(0) 
                           => n_1107);
   muxi_3 : MUX51_GENERIC_NBIT16_1 port map( A0(15) => set_signal_3_1_15_port, 
                           A0(14) => set_signal_3_1_14_port, A0(13) => 
                           set_signal_3_1_13_port, A0(12) => 
                           set_signal_3_1_12_port, A0(11) => 
                           set_signal_3_1_11_port, A0(10) => 
                           set_signal_3_1_10_port, A0(9) => 
                           set_signal_3_1_9_port, A0(8) => 
                           set_signal_3_1_8_port, A0(7) => 
                           set_signal_3_1_7_port, A0(6) => 
                           set_signal_3_1_6_port, A0(5) => 
                           set_signal_3_1_5_port, A0(4) => 
                           set_signal_3_1_4_port, A0(3) => 
                           set_signal_3_1_3_port, A0(2) => 
                           set_signal_3_1_2_port, A0(1) => 
                           set_signal_3_1_1_port, A0(0) => 
                           set_signal_3_1_0_port, A1(15) => 
                           set_signal_3_2_15_port, A1(14) => 
                           set_signal_3_2_14_port, A1(13) => 
                           set_signal_3_2_13_port, A1(12) => 
                           set_signal_3_2_12_port, A1(11) => 
                           set_signal_3_2_11_port, A1(10) => 
                           set_signal_3_2_10_port, A1(9) => 
                           set_signal_3_2_9_port, A1(8) => 
                           set_signal_3_2_8_port, A1(7) => 
                           set_signal_3_2_7_port, A1(6) => 
                           set_signal_3_2_6_port, A1(5) => 
                           set_signal_3_2_5_port, A1(4) => 
                           set_signal_3_2_4_port, A1(3) => 
                           set_signal_3_2_3_port, A1(2) => 
                           set_signal_3_2_2_port, A1(1) => 
                           set_signal_3_2_1_port, A1(0) => 
                           set_signal_3_2_0_port, A2(15) => 
                           set_signal_3_3_15_port, A2(14) => 
                           set_signal_3_3_14_port, A2(13) => 
                           set_signal_3_3_13_port, A2(12) => 
                           set_signal_3_3_12_port, A2(11) => 
                           set_signal_3_3_11_port, A2(10) => 
                           set_signal_3_3_10_port, A2(9) => 
                           set_signal_3_3_9_port, A2(8) => 
                           set_signal_3_3_8_port, A2(7) => 
                           set_signal_3_3_7_port, A2(6) => 
                           set_signal_3_3_6_port, A2(5) => 
                           set_signal_3_3_5_port, A2(4) => 
                           set_signal_3_3_4_port, A2(3) => 
                           set_signal_3_3_3_port, A2(2) => 
                           set_signal_3_3_2_port, A2(1) => 
                           set_signal_3_3_1_port, A2(0) => 
                           set_signal_3_3_0_port, A3(15) => 
                           set_signal_3_4_15_port, A3(14) => 
                           set_signal_3_4_14_port, A3(13) => 
                           set_signal_3_4_13_port, A3(12) => 
                           set_signal_3_4_12_port, A3(11) => 
                           set_signal_3_4_11_port, A3(10) => 
                           set_signal_3_4_10_port, A3(9) => 
                           set_signal_3_4_9_port, A3(8) => 
                           set_signal_3_4_8_port, A3(7) => 
                           set_signal_3_4_7_port, A3(6) => 
                           set_signal_3_4_6_port, A3(5) => 
                           set_signal_3_4_5_port, A3(4) => 
                           set_signal_3_4_4_port, A3(3) => 
                           set_signal_3_4_3_port, A3(2) => 
                           set_signal_3_4_2_port, A3(1) => 
                           set_signal_3_4_1_port, A3(0) => 
                           set_signal_3_4_0_port, A4(15) => 
                           set_signal_3_5_15_port, A4(14) => 
                           set_signal_3_5_14_port, A4(13) => 
                           set_signal_3_5_13_port, A4(12) => 
                           set_signal_3_5_12_port, A4(11) => 
                           set_signal_3_5_11_port, A4(10) => 
                           set_signal_3_5_10_port, A4(9) => 
                           set_signal_3_5_9_port, A4(8) => 
                           set_signal_3_5_8_port, A4(7) => 
                           set_signal_3_5_7_port, A4(6) => 
                           set_signal_3_5_6_port, A4(5) => 
                           set_signal_3_5_5_port, A4(4) => 
                           set_signal_3_5_4_port, A4(3) => 
                           set_signal_3_5_3_port, A4(2) => 
                           set_signal_3_5_2_port, A4(1) => 
                           set_signal_3_5_1_port, A4(0) => 
                           set_signal_3_5_0_port, SEL(2) => 
                           enc_signal_3_1_2_port, SEL(1) => 
                           enc_signal_3_1_1_port, SEL(0) => 
                           enc_signal_3_1_0_port, Y(15) => 
                           rca_signal_3_0_15_port, Y(14) => 
                           rca_signal_3_0_14_port, Y(13) => 
                           rca_signal_3_0_13_port, Y(12) => 
                           rca_signal_3_0_12_port, Y(11) => 
                           rca_signal_3_0_11_port, Y(10) => 
                           rca_signal_3_0_10_port, Y(9) => 
                           rca_signal_3_0_9_port, Y(8) => rca_signal_3_0_8_port
                           , Y(7) => rca_signal_3_0_7_port, Y(6) => 
                           rca_signal_3_0_6_port, Y(5) => rca_signal_3_0_5_port
                           , Y(4) => rca_signal_3_0_4_port, Y(3) => 
                           rca_signal_3_0_3_port, Y(2) => rca_signal_3_0_2_port
                           , Y(1) => rca_signal_3_0_1_port, Y(0) => 
                           rca_signal_3_0_0_port);
   rcai_3 : RCA_size16_1 port map( a(15) => rca_signal_3_0_15_port, a(14) => 
                           rca_signal_3_0_14_port, a(13) => 
                           rca_signal_3_0_13_port, a(12) => 
                           rca_signal_3_0_12_port, a(11) => 
                           rca_signal_3_0_11_port, a(10) => 
                           rca_signal_3_0_10_port, a(9) => 
                           rca_signal_3_0_9_port, a(8) => rca_signal_3_0_8_port
                           , a(7) => rca_signal_3_0_7_port, a(6) => 
                           rca_signal_3_0_6_port, a(5) => rca_signal_3_0_5_port
                           , a(4) => rca_signal_3_0_4_port, a(3) => 
                           rca_signal_3_0_3_port, a(2) => rca_signal_3_0_2_port
                           , a(1) => rca_signal_3_0_1_port, a(0) => 
                           rca_signal_3_0_0_port, b(15) => 
                           rca_signal_3_1_15_port, b(14) => 
                           rca_signal_3_1_14_port, b(13) => 
                           rca_signal_3_1_13_port, b(12) => 
                           rca_signal_3_1_12_port, b(11) => 
                           rca_signal_3_1_11_port, b(10) => 
                           rca_signal_3_1_10_port, b(9) => 
                           rca_signal_3_1_9_port, b(8) => rca_signal_3_1_8_port
                           , b(7) => rca_signal_3_1_7_port, b(6) => 
                           rca_signal_3_1_6_port, b(5) => rca_signal_3_1_5_port
                           , b(4) => rca_signal_3_1_4_port, b(3) => 
                           rca_signal_3_1_3_port, b(2) => rca_signal_3_1_2_port
                           , b(1) => rca_signal_3_1_1_port, b(0) => 
                           rca_signal_3_1_0_port, c_in => X_Logic0_port, c_out 
                           => n_1108, sum(15) => Y_mp(15), sum(14) => Y_mp(14),
                           sum(13) => Y_mp(13), sum(12) => Y_mp(12), sum(11) =>
                           Y_mp(11), sum(10) => Y_mp(10), sum(9) => Y_mp(9), 
                           sum(8) => Y_mp(8), sum(7) => Y_mp(7), sum(6) => 
                           Y_mp(6), sum(5) => Y_mp(5), sum(4) => Y_mp(4), 
                           sum(3) => Y_mp(3), sum(2) => Y_mp(2), sum(1) => 
                           Y_mp(1), sum(0) => Y_mp(0));
   set_signal_1_6_0_port <= '0';
   set_signal_1_6_1_port <= '0';
   set_signal_1_5_0_port <= '0';
   set_signal_1_4_0_port <= '0';
   set_signal_1_1_0_port <= '0';
   set_signal_1_1_1_port <= '0';
   set_signal_1_1_2_port <= '0';
   set_signal_1_1_3_port <= '0';
   set_signal_1_1_4_port <= '0';
   set_signal_1_1_5_port <= '0';
   set_signal_1_1_6_port <= '0';
   set_signal_1_1_7_port <= '0';
   set_signal_1_1_8_port <= '0';
   set_signal_1_1_9_port <= '0';
   set_signal_1_1_10_port <= '0';
   set_signal_1_1_11_port <= '0';
   set_signal_1_1_12_port <= '0';
   set_signal_1_1_13_port <= '0';
   set_signal_1_1_14_port <= '0';
   set_signal_1_1_15_port <= '0';
   set_signal_2_6_0_port <= '0';
   set_signal_2_6_1_port <= '0';
   set_signal_2_5_0_port <= '0';
   set_signal_2_4_0_port <= '0';
   set_signal_2_1_0_port <= '0';
   set_signal_2_1_1_port <= '0';
   set_signal_2_1_2_port <= '0';
   set_signal_2_1_3_port <= '0';
   set_signal_2_1_4_port <= '0';
   set_signal_2_1_5_port <= '0';
   set_signal_2_1_6_port <= '0';
   set_signal_2_1_7_port <= '0';
   set_signal_2_1_8_port <= '0';
   set_signal_2_1_9_port <= '0';
   set_signal_2_1_10_port <= '0';
   set_signal_2_1_11_port <= '0';
   set_signal_2_1_12_port <= '0';
   set_signal_2_1_13_port <= '0';
   set_signal_2_1_14_port <= '0';
   set_signal_2_1_15_port <= '0';
   set_signal_3_5_0_port <= '0';
   set_signal_3_4_0_port <= '0';
   set_signal_3_1_0_port <= '0';
   set_signal_3_1_1_port <= '0';
   set_signal_3_1_2_port <= '0';
   set_signal_3_1_3_port <= '0';
   set_signal_3_1_4_port <= '0';
   set_signal_3_1_5_port <= '0';
   set_signal_3_1_6_port <= '0';
   set_signal_3_1_7_port <= '0';
   set_signal_3_1_8_port <= '0';
   set_signal_3_1_9_port <= '0';
   set_signal_3_1_10_port <= '0';
   set_signal_3_1_11_port <= '0';
   set_signal_3_1_12_port <= '0';
   set_signal_3_1_13_port <= '0';
   set_signal_3_1_14_port <= '0';
   set_signal_3_1_15_port <= '0';
   set_signal_0_6_0_port <= '0';
   set_signal_0_6_1_port <= '0';
   set_signal_0_5_0_port <= '0';
   set_signal_0_4_0_port <= '0';
   set_signal_0_1_0_port <= '0';
   set_signal_0_1_1_port <= '0';
   set_signal_0_1_2_port <= '0';
   set_signal_0_1_3_port <= '0';
   set_signal_0_1_4_port <= '0';
   set_signal_0_1_5_port <= '0';
   set_signal_0_1_6_port <= '0';
   set_signal_0_1_7_port <= '0';
   set_signal_0_1_8_port <= '0';
   set_signal_0_1_9_port <= '0';
   set_signal_0_1_10_port <= '0';
   set_signal_0_1_11_port <= '0';
   set_signal_0_1_12_port <= '0';
   set_signal_0_1_13_port <= '0';
   set_signal_0_1_14_port <= '0';
   set_signal_0_1_15_port <= '0';

end SYN_STRUCTURAL;
