
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_topLevel_1 is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_topLevel_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_topLevel_1.all;

entity register_file_WORD_SIZE32_ADDR_SIZE6 is

   port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
         ADD_RD2 : in std_logic_vector (5 downto 0);  DATAIN : in 
         std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector (31
         downto 0));

end register_file_WORD_SIZE32_ADDR_SIZE6;

architecture SYN_Beh of register_file_WORD_SIZE32_ADDR_SIZE6 is

   component GTECH_NOT
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component GTECH_AND2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component SELECT_OP
      generic( num_inputs, input_width : integer );
      port( DATA : in std_logic_vector( num_inputs* input_width - 1 downto 0 );
            CONTROL : in std_logic_vector( num_inputs - 1 downto 0 ); Z : out 
            std_logic_vector( input_width - 1 downto 0 ) );
   end component;
   
   component GTECH_BUF
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
      generic ( ac_as_q, ac_as_qn, sc_ss_q : integer );
      port(
         clear, preset, enable, data_in, synch_clear, synch_preset, 
            synch_toggle, synch_enable, next_state, clocked_on : in std_logic;
         Q, QN : buffer std_logic
      );
   end component;
   
   signal N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
      X_Logic1_port, X_Logic0_port, CLK_port, RD1_port, RD2_port, 
      DATAIN_31_port, DATAIN_30_port, DATAIN_29_port, DATAIN_28_port, 
      DATAIN_27_port, DATAIN_26_port, DATAIN_25_port, DATAIN_24_port, 
      DATAIN_23_port, DATAIN_22_port, DATAIN_21_port, DATAIN_20_port, 
      DATAIN_19_port, DATAIN_18_port, DATAIN_17_port, DATAIN_16_port, 
      DATAIN_15_port, DATAIN_14_port, DATAIN_13_port, DATAIN_12_port, 
      DATAIN_11_port, DATAIN_10_port, DATAIN_9_port, DATAIN_8_port, 
      DATAIN_7_port, DATAIN_6_port, DATAIN_5_port, DATAIN_4_port, DATAIN_3_port
      , DATAIN_2_port, DATAIN_1_port, DATAIN_0_port, OUT1_31_port, OUT1_30_port
      , OUT1_29_port, OUT1_28_port, OUT1_27_port, OUT1_26_port, OUT1_25_port, 
      OUT1_24_port, OUT1_23_port, OUT1_22_port, OUT1_21_port, OUT1_20_port, 
      OUT1_19_port, OUT1_18_port, OUT1_17_port, OUT1_16_port, OUT1_15_port, 
      OUT1_14_port, OUT1_13_port, OUT1_12_port, OUT1_11_port, OUT1_10_port, 
      OUT1_9_port, OUT1_8_port, OUT1_7_port, OUT1_6_port, OUT1_5_port, 
      OUT1_4_port, OUT1_3_port, OUT1_2_port, OUT1_1_port, OUT1_0_port, 
      OUT2_31_port, OUT2_30_port, OUT2_29_port, OUT2_28_port, OUT2_27_port, 
      OUT2_26_port, OUT2_25_port, OUT2_24_port, OUT2_23_port, OUT2_22_port, 
      OUT2_21_port, OUT2_20_port, OUT2_19_port, OUT2_18_port, OUT2_17_port, 
      OUT2_16_port, OUT2_15_port, OUT2_14_port, OUT2_13_port, OUT2_12_port, 
      OUT2_11_port, OUT2_10_port, OUT2_9_port, OUT2_8_port, OUT2_7_port, 
      OUT2_6_port, OUT2_5_port, OUT2_4_port, OUT2_3_port, OUT2_2_port, 
      OUT2_1_port, OUT2_0_port, N16, REGISTERS_0_31_port, REGISTERS_0_30_port, 
      REGISTERS_0_29_port, REGISTERS_0_28_port, REGISTERS_0_27_port, 
      REGISTERS_0_26_port, REGISTERS_0_25_port, REGISTERS_0_24_port, 
      REGISTERS_0_23_port, REGISTERS_0_22_port, REGISTERS_0_21_port, 
      REGISTERS_0_20_port, REGISTERS_0_19_port, REGISTERS_0_18_port, 
      REGISTERS_0_17_port, REGISTERS_0_16_port, REGISTERS_0_15_port, 
      REGISTERS_0_14_port, REGISTERS_0_13_port, REGISTERS_0_12_port, 
      REGISTERS_0_11_port, REGISTERS_0_10_port, REGISTERS_0_9_port, 
      REGISTERS_0_8_port, REGISTERS_0_7_port, REGISTERS_0_6_port, 
      REGISTERS_0_5_port, REGISTERS_0_4_port, REGISTERS_0_3_port, 
      REGISTERS_0_2_port, REGISTERS_0_1_port, REGISTERS_0_0_port, 
      REGISTERS_1_31_port, REGISTERS_1_30_port, REGISTERS_1_29_port, 
      REGISTERS_1_28_port, REGISTERS_1_27_port, REGISTERS_1_26_port, 
      REGISTERS_1_25_port, REGISTERS_1_24_port, REGISTERS_1_23_port, 
      REGISTERS_1_22_port, REGISTERS_1_21_port, REGISTERS_1_20_port, 
      REGISTERS_1_19_port, REGISTERS_1_18_port, REGISTERS_1_17_port, 
      REGISTERS_1_16_port, REGISTERS_1_15_port, REGISTERS_1_14_port, 
      REGISTERS_1_13_port, REGISTERS_1_12_port, REGISTERS_1_11_port, 
      REGISTERS_1_10_port, REGISTERS_1_9_port, REGISTERS_1_8_port, 
      REGISTERS_1_7_port, REGISTERS_1_6_port, REGISTERS_1_5_port, 
      REGISTERS_1_4_port, REGISTERS_1_3_port, REGISTERS_1_2_port, 
      REGISTERS_1_1_port, REGISTERS_1_0_port, REGISTERS_2_31_port, 
      REGISTERS_2_30_port, REGISTERS_2_29_port, REGISTERS_2_28_port, 
      REGISTERS_2_27_port, REGISTERS_2_26_port, REGISTERS_2_25_port, 
      REGISTERS_2_24_port, REGISTERS_2_23_port, REGISTERS_2_22_port, 
      REGISTERS_2_21_port, REGISTERS_2_20_port, REGISTERS_2_19_port, 
      REGISTERS_2_18_port, REGISTERS_2_17_port, REGISTERS_2_16_port, 
      REGISTERS_2_15_port, REGISTERS_2_14_port, REGISTERS_2_13_port, 
      REGISTERS_2_12_port, REGISTERS_2_11_port, REGISTERS_2_10_port, 
      REGISTERS_2_9_port, REGISTERS_2_8_port, REGISTERS_2_7_port, 
      REGISTERS_2_6_port, REGISTERS_2_5_port, REGISTERS_2_4_port, 
      REGISTERS_2_3_port, REGISTERS_2_2_port, REGISTERS_2_1_port, 
      REGISTERS_2_0_port, REGISTERS_3_31_port, REGISTERS_3_30_port, 
      REGISTERS_3_29_port, REGISTERS_3_28_port, REGISTERS_3_27_port, 
      REGISTERS_3_26_port, REGISTERS_3_25_port, REGISTERS_3_24_port, 
      REGISTERS_3_23_port, REGISTERS_3_22_port, REGISTERS_3_21_port, 
      REGISTERS_3_20_port, REGISTERS_3_19_port, REGISTERS_3_18_port, 
      REGISTERS_3_17_port, REGISTERS_3_16_port, REGISTERS_3_15_port, 
      REGISTERS_3_14_port, REGISTERS_3_13_port, REGISTERS_3_12_port, 
      REGISTERS_3_11_port, REGISTERS_3_10_port, REGISTERS_3_9_port, 
      REGISTERS_3_8_port, REGISTERS_3_7_port, REGISTERS_3_6_port, 
      REGISTERS_3_5_port, REGISTERS_3_4_port, REGISTERS_3_3_port, 
      REGISTERS_3_2_port, REGISTERS_3_1_port, REGISTERS_3_0_port, 
      REGISTERS_4_31_port, REGISTERS_4_30_port, REGISTERS_4_29_port, 
      REGISTERS_4_28_port, REGISTERS_4_27_port, REGISTERS_4_26_port, 
      REGISTERS_4_25_port, REGISTERS_4_24_port, REGISTERS_4_23_port, 
      REGISTERS_4_22_port, REGISTERS_4_21_port, REGISTERS_4_20_port, 
      REGISTERS_4_19_port, REGISTERS_4_18_port, REGISTERS_4_17_port, 
      REGISTERS_4_16_port, REGISTERS_4_15_port, REGISTERS_4_14_port, 
      REGISTERS_4_13_port, REGISTERS_4_12_port, REGISTERS_4_11_port, 
      REGISTERS_4_10_port, REGISTERS_4_9_port, REGISTERS_4_8_port, 
      REGISTERS_4_7_port, REGISTERS_4_6_port, REGISTERS_4_5_port, 
      REGISTERS_4_4_port, REGISTERS_4_3_port, REGISTERS_4_2_port, 
      REGISTERS_4_1_port, REGISTERS_4_0_port, REGISTERS_5_31_port, 
      REGISTERS_5_30_port, REGISTERS_5_29_port, REGISTERS_5_28_port, 
      REGISTERS_5_27_port, REGISTERS_5_26_port, REGISTERS_5_25_port, 
      REGISTERS_5_24_port, REGISTERS_5_23_port, REGISTERS_5_22_port, 
      REGISTERS_5_21_port, REGISTERS_5_20_port, REGISTERS_5_19_port, 
      REGISTERS_5_18_port, REGISTERS_5_17_port, REGISTERS_5_16_port, 
      REGISTERS_5_15_port, REGISTERS_5_14_port, REGISTERS_5_13_port, 
      REGISTERS_5_12_port, REGISTERS_5_11_port, REGISTERS_5_10_port, 
      REGISTERS_5_9_port, REGISTERS_5_8_port, REGISTERS_5_7_port, 
      REGISTERS_5_6_port, REGISTERS_5_5_port, REGISTERS_5_4_port, 
      REGISTERS_5_3_port, REGISTERS_5_2_port, REGISTERS_5_1_port, 
      REGISTERS_5_0_port, REGISTERS_6_31_port, REGISTERS_6_30_port, 
      REGISTERS_6_29_port, REGISTERS_6_28_port, REGISTERS_6_27_port, 
      REGISTERS_6_26_port, REGISTERS_6_25_port, REGISTERS_6_24_port, 
      REGISTERS_6_23_port, REGISTERS_6_22_port, REGISTERS_6_21_port, 
      REGISTERS_6_20_port, REGISTERS_6_19_port, REGISTERS_6_18_port, 
      REGISTERS_6_17_port, REGISTERS_6_16_port, REGISTERS_6_15_port, 
      REGISTERS_6_14_port, REGISTERS_6_13_port, REGISTERS_6_12_port, 
      REGISTERS_6_11_port, REGISTERS_6_10_port, REGISTERS_6_9_port, 
      REGISTERS_6_8_port, REGISTERS_6_7_port, REGISTERS_6_6_port, 
      REGISTERS_6_5_port, REGISTERS_6_4_port, REGISTERS_6_3_port, 
      REGISTERS_6_2_port, REGISTERS_6_1_port, REGISTERS_6_0_port, 
      REGISTERS_7_31_port, REGISTERS_7_30_port, REGISTERS_7_29_port, 
      REGISTERS_7_28_port, REGISTERS_7_27_port, REGISTERS_7_26_port, 
      REGISTERS_7_25_port, REGISTERS_7_24_port, REGISTERS_7_23_port, 
      REGISTERS_7_22_port, REGISTERS_7_21_port, REGISTERS_7_20_port, 
      REGISTERS_7_19_port, REGISTERS_7_18_port, REGISTERS_7_17_port, 
      REGISTERS_7_16_port, REGISTERS_7_15_port, REGISTERS_7_14_port, 
      REGISTERS_7_13_port, REGISTERS_7_12_port, REGISTERS_7_11_port, 
      REGISTERS_7_10_port, REGISTERS_7_9_port, REGISTERS_7_8_port, 
      REGISTERS_7_7_port, REGISTERS_7_6_port, REGISTERS_7_5_port, 
      REGISTERS_7_4_port, REGISTERS_7_3_port, REGISTERS_7_2_port, 
      REGISTERS_7_1_port, REGISTERS_7_0_port, REGISTERS_8_31_port, 
      REGISTERS_8_30_port, REGISTERS_8_29_port, REGISTERS_8_28_port, 
      REGISTERS_8_27_port, REGISTERS_8_26_port, REGISTERS_8_25_port, 
      REGISTERS_8_24_port, REGISTERS_8_23_port, REGISTERS_8_22_port, 
      REGISTERS_8_21_port, REGISTERS_8_20_port, REGISTERS_8_19_port, 
      REGISTERS_8_18_port, REGISTERS_8_17_port, REGISTERS_8_16_port, 
      REGISTERS_8_15_port, REGISTERS_8_14_port, REGISTERS_8_13_port, 
      REGISTERS_8_12_port, REGISTERS_8_11_port, REGISTERS_8_10_port, 
      REGISTERS_8_9_port, REGISTERS_8_8_port, REGISTERS_8_7_port, 
      REGISTERS_8_6_port, REGISTERS_8_5_port, REGISTERS_8_4_port, 
      REGISTERS_8_3_port, REGISTERS_8_2_port, REGISTERS_8_1_port, 
      REGISTERS_8_0_port, REGISTERS_9_31_port, REGISTERS_9_30_port, 
      REGISTERS_9_29_port, REGISTERS_9_28_port, REGISTERS_9_27_port, 
      REGISTERS_9_26_port, REGISTERS_9_25_port, REGISTERS_9_24_port, 
      REGISTERS_9_23_port, REGISTERS_9_22_port, REGISTERS_9_21_port, 
      REGISTERS_9_20_port, REGISTERS_9_19_port, REGISTERS_9_18_port, 
      REGISTERS_9_17_port, REGISTERS_9_16_port, REGISTERS_9_15_port, 
      REGISTERS_9_14_port, REGISTERS_9_13_port, REGISTERS_9_12_port, 
      REGISTERS_9_11_port, REGISTERS_9_10_port, REGISTERS_9_9_port, 
      REGISTERS_9_8_port, REGISTERS_9_7_port, REGISTERS_9_6_port, 
      REGISTERS_9_5_port, REGISTERS_9_4_port, REGISTERS_9_3_port, 
      REGISTERS_9_2_port, REGISTERS_9_1_port, REGISTERS_9_0_port, 
      REGISTERS_10_31_port, REGISTERS_10_30_port, REGISTERS_10_29_port, 
      REGISTERS_10_28_port, REGISTERS_10_27_port, REGISTERS_10_26_port, 
      REGISTERS_10_25_port, REGISTERS_10_24_port, REGISTERS_10_23_port, 
      REGISTERS_10_22_port, REGISTERS_10_21_port, REGISTERS_10_20_port, 
      REGISTERS_10_19_port, REGISTERS_10_18_port, REGISTERS_10_17_port, 
      REGISTERS_10_16_port, REGISTERS_10_15_port, REGISTERS_10_14_port, 
      REGISTERS_10_13_port, REGISTERS_10_12_port, REGISTERS_10_11_port, 
      REGISTERS_10_10_port, REGISTERS_10_9_port, REGISTERS_10_8_port, 
      REGISTERS_10_7_port, REGISTERS_10_6_port, REGISTERS_10_5_port, 
      REGISTERS_10_4_port, REGISTERS_10_3_port, REGISTERS_10_2_port, 
      REGISTERS_10_1_port, REGISTERS_10_0_port, REGISTERS_11_31_port, 
      REGISTERS_11_30_port, REGISTERS_11_29_port, REGISTERS_11_28_port, 
      REGISTERS_11_27_port, REGISTERS_11_26_port, REGISTERS_11_25_port, 
      REGISTERS_11_24_port, REGISTERS_11_23_port, REGISTERS_11_22_port, 
      REGISTERS_11_21_port, REGISTERS_11_20_port, REGISTERS_11_19_port, 
      REGISTERS_11_18_port, REGISTERS_11_17_port, REGISTERS_11_16_port, 
      REGISTERS_11_15_port, REGISTERS_11_14_port, REGISTERS_11_13_port, 
      REGISTERS_11_12_port, REGISTERS_11_11_port, REGISTERS_11_10_port, 
      REGISTERS_11_9_port, REGISTERS_11_8_port, REGISTERS_11_7_port, 
      REGISTERS_11_6_port, REGISTERS_11_5_port, REGISTERS_11_4_port, 
      REGISTERS_11_3_port, REGISTERS_11_2_port, REGISTERS_11_1_port, 
      REGISTERS_11_0_port, REGISTERS_12_31_port, REGISTERS_12_30_port, 
      REGISTERS_12_29_port, REGISTERS_12_28_port, REGISTERS_12_27_port, 
      REGISTERS_12_26_port, REGISTERS_12_25_port, REGISTERS_12_24_port, 
      REGISTERS_12_23_port, REGISTERS_12_22_port, REGISTERS_12_21_port, 
      REGISTERS_12_20_port, REGISTERS_12_19_port, REGISTERS_12_18_port, 
      REGISTERS_12_17_port, REGISTERS_12_16_port, REGISTERS_12_15_port, 
      REGISTERS_12_14_port, REGISTERS_12_13_port, REGISTERS_12_12_port, 
      REGISTERS_12_11_port, REGISTERS_12_10_port, REGISTERS_12_9_port, 
      REGISTERS_12_8_port, REGISTERS_12_7_port, REGISTERS_12_6_port, 
      REGISTERS_12_5_port, REGISTERS_12_4_port, REGISTERS_12_3_port, 
      REGISTERS_12_2_port, REGISTERS_12_1_port, REGISTERS_12_0_port, 
      REGISTERS_13_31_port, REGISTERS_13_30_port, REGISTERS_13_29_port, 
      REGISTERS_13_28_port, REGISTERS_13_27_port, REGISTERS_13_26_port, 
      REGISTERS_13_25_port, REGISTERS_13_24_port, REGISTERS_13_23_port, 
      REGISTERS_13_22_port, REGISTERS_13_21_port, REGISTERS_13_20_port, 
      REGISTERS_13_19_port, REGISTERS_13_18_port, REGISTERS_13_17_port, 
      REGISTERS_13_16_port, REGISTERS_13_15_port, REGISTERS_13_14_port, 
      REGISTERS_13_13_port, REGISTERS_13_12_port, REGISTERS_13_11_port, 
      REGISTERS_13_10_port, REGISTERS_13_9_port, REGISTERS_13_8_port, 
      REGISTERS_13_7_port, REGISTERS_13_6_port, REGISTERS_13_5_port, 
      REGISTERS_13_4_port, REGISTERS_13_3_port, REGISTERS_13_2_port, 
      REGISTERS_13_1_port, REGISTERS_13_0_port, REGISTERS_14_31_port, 
      REGISTERS_14_30_port, REGISTERS_14_29_port, REGISTERS_14_28_port, 
      REGISTERS_14_27_port, REGISTERS_14_26_port, REGISTERS_14_25_port, 
      REGISTERS_14_24_port, REGISTERS_14_23_port, REGISTERS_14_22_port, 
      REGISTERS_14_21_port, REGISTERS_14_20_port, REGISTERS_14_19_port, 
      REGISTERS_14_18_port, REGISTERS_14_17_port, REGISTERS_14_16_port, 
      REGISTERS_14_15_port, REGISTERS_14_14_port, REGISTERS_14_13_port, 
      REGISTERS_14_12_port, REGISTERS_14_11_port, REGISTERS_14_10_port, 
      REGISTERS_14_9_port, REGISTERS_14_8_port, REGISTERS_14_7_port, 
      REGISTERS_14_6_port, REGISTERS_14_5_port, REGISTERS_14_4_port, 
      REGISTERS_14_3_port, REGISTERS_14_2_port, REGISTERS_14_1_port, 
      REGISTERS_14_0_port, REGISTERS_15_31_port, REGISTERS_15_30_port, 
      REGISTERS_15_29_port, REGISTERS_15_28_port, REGISTERS_15_27_port, 
      REGISTERS_15_26_port, REGISTERS_15_25_port, REGISTERS_15_24_port, 
      REGISTERS_15_23_port, REGISTERS_15_22_port, REGISTERS_15_21_port, 
      REGISTERS_15_20_port, REGISTERS_15_19_port, REGISTERS_15_18_port, 
      REGISTERS_15_17_port, REGISTERS_15_16_port, REGISTERS_15_15_port, 
      REGISTERS_15_14_port, REGISTERS_15_13_port, REGISTERS_15_12_port, 
      REGISTERS_15_11_port, REGISTERS_15_10_port, REGISTERS_15_9_port, 
      REGISTERS_15_8_port, REGISTERS_15_7_port, REGISTERS_15_6_port, 
      REGISTERS_15_5_port, REGISTERS_15_4_port, REGISTERS_15_3_port, 
      REGISTERS_15_2_port, REGISTERS_15_1_port, REGISTERS_15_0_port, 
      REGISTERS_16_31_port, REGISTERS_16_30_port, REGISTERS_16_29_port, 
      REGISTERS_16_28_port, REGISTERS_16_27_port, REGISTERS_16_26_port, 
      REGISTERS_16_25_port, REGISTERS_16_24_port, REGISTERS_16_23_port, 
      REGISTERS_16_22_port, REGISTERS_16_21_port, REGISTERS_16_20_port, 
      REGISTERS_16_19_port, REGISTERS_16_18_port, REGISTERS_16_17_port, 
      REGISTERS_16_16_port, REGISTERS_16_15_port, REGISTERS_16_14_port, 
      REGISTERS_16_13_port, REGISTERS_16_12_port, REGISTERS_16_11_port, 
      REGISTERS_16_10_port, REGISTERS_16_9_port, REGISTERS_16_8_port, 
      REGISTERS_16_7_port, REGISTERS_16_6_port, REGISTERS_16_5_port, 
      REGISTERS_16_4_port, REGISTERS_16_3_port, REGISTERS_16_2_port, 
      REGISTERS_16_1_port, REGISTERS_16_0_port, REGISTERS_17_31_port, 
      REGISTERS_17_30_port, REGISTERS_17_29_port, REGISTERS_17_28_port, 
      REGISTERS_17_27_port, REGISTERS_17_26_port, REGISTERS_17_25_port, 
      REGISTERS_17_24_port, REGISTERS_17_23_port, REGISTERS_17_22_port, 
      REGISTERS_17_21_port, REGISTERS_17_20_port, REGISTERS_17_19_port, 
      REGISTERS_17_18_port, REGISTERS_17_17_port, REGISTERS_17_16_port, 
      REGISTERS_17_15_port, REGISTERS_17_14_port, REGISTERS_17_13_port, 
      REGISTERS_17_12_port, REGISTERS_17_11_port, REGISTERS_17_10_port, 
      REGISTERS_17_9_port, REGISTERS_17_8_port, REGISTERS_17_7_port, 
      REGISTERS_17_6_port, REGISTERS_17_5_port, REGISTERS_17_4_port, 
      REGISTERS_17_3_port, REGISTERS_17_2_port, REGISTERS_17_1_port, 
      REGISTERS_17_0_port, REGISTERS_18_31_port, REGISTERS_18_30_port, 
      REGISTERS_18_29_port, REGISTERS_18_28_port, REGISTERS_18_27_port, 
      REGISTERS_18_26_port, REGISTERS_18_25_port, REGISTERS_18_24_port, 
      REGISTERS_18_23_port, REGISTERS_18_22_port, REGISTERS_18_21_port, 
      REGISTERS_18_20_port, REGISTERS_18_19_port, REGISTERS_18_18_port, 
      REGISTERS_18_17_port, REGISTERS_18_16_port, REGISTERS_18_15_port, 
      REGISTERS_18_14_port, REGISTERS_18_13_port, REGISTERS_18_12_port, 
      REGISTERS_18_11_port, REGISTERS_18_10_port, REGISTERS_18_9_port, 
      REGISTERS_18_8_port, REGISTERS_18_7_port, REGISTERS_18_6_port, 
      REGISTERS_18_5_port, REGISTERS_18_4_port, REGISTERS_18_3_port, 
      REGISTERS_18_2_port, REGISTERS_18_1_port, REGISTERS_18_0_port, 
      REGISTERS_19_31_port, REGISTERS_19_30_port, REGISTERS_19_29_port, 
      REGISTERS_19_28_port, REGISTERS_19_27_port, REGISTERS_19_26_port, 
      REGISTERS_19_25_port, REGISTERS_19_24_port, REGISTERS_19_23_port, 
      REGISTERS_19_22_port, REGISTERS_19_21_port, REGISTERS_19_20_port, 
      REGISTERS_19_19_port, REGISTERS_19_18_port, REGISTERS_19_17_port, 
      REGISTERS_19_16_port, REGISTERS_19_15_port, REGISTERS_19_14_port, 
      REGISTERS_19_13_port, REGISTERS_19_12_port, REGISTERS_19_11_port, 
      REGISTERS_19_10_port, REGISTERS_19_9_port, REGISTERS_19_8_port, 
      REGISTERS_19_7_port, REGISTERS_19_6_port, REGISTERS_19_5_port, 
      REGISTERS_19_4_port, REGISTERS_19_3_port, REGISTERS_19_2_port, 
      REGISTERS_19_1_port, REGISTERS_19_0_port, REGISTERS_20_31_port, 
      REGISTERS_20_30_port, REGISTERS_20_29_port, REGISTERS_20_28_port, 
      REGISTERS_20_27_port, REGISTERS_20_26_port, REGISTERS_20_25_port, 
      REGISTERS_20_24_port, REGISTERS_20_23_port, REGISTERS_20_22_port, 
      REGISTERS_20_21_port, REGISTERS_20_20_port, REGISTERS_20_19_port, 
      REGISTERS_20_18_port, REGISTERS_20_17_port, REGISTERS_20_16_port, 
      REGISTERS_20_15_port, REGISTERS_20_14_port, REGISTERS_20_13_port, 
      REGISTERS_20_12_port, REGISTERS_20_11_port, REGISTERS_20_10_port, 
      REGISTERS_20_9_port, REGISTERS_20_8_port, REGISTERS_20_7_port, 
      REGISTERS_20_6_port, REGISTERS_20_5_port, REGISTERS_20_4_port, 
      REGISTERS_20_3_port, REGISTERS_20_2_port, REGISTERS_20_1_port, 
      REGISTERS_20_0_port, REGISTERS_21_31_port, REGISTERS_21_30_port, 
      REGISTERS_21_29_port, REGISTERS_21_28_port, REGISTERS_21_27_port, 
      REGISTERS_21_26_port, REGISTERS_21_25_port, REGISTERS_21_24_port, 
      REGISTERS_21_23_port, REGISTERS_21_22_port, REGISTERS_21_21_port, 
      REGISTERS_21_20_port, REGISTERS_21_19_port, REGISTERS_21_18_port, 
      REGISTERS_21_17_port, REGISTERS_21_16_port, REGISTERS_21_15_port, 
      REGISTERS_21_14_port, REGISTERS_21_13_port, REGISTERS_21_12_port, 
      REGISTERS_21_11_port, REGISTERS_21_10_port, REGISTERS_21_9_port, 
      REGISTERS_21_8_port, REGISTERS_21_7_port, REGISTERS_21_6_port, 
      REGISTERS_21_5_port, REGISTERS_21_4_port, REGISTERS_21_3_port, 
      REGISTERS_21_2_port, REGISTERS_21_1_port, REGISTERS_21_0_port, 
      REGISTERS_22_31_port, REGISTERS_22_30_port, REGISTERS_22_29_port, 
      REGISTERS_22_28_port, REGISTERS_22_27_port, REGISTERS_22_26_port, 
      REGISTERS_22_25_port, REGISTERS_22_24_port, REGISTERS_22_23_port, 
      REGISTERS_22_22_port, REGISTERS_22_21_port, REGISTERS_22_20_port, 
      REGISTERS_22_19_port, REGISTERS_22_18_port, REGISTERS_22_17_port, 
      REGISTERS_22_16_port, REGISTERS_22_15_port, REGISTERS_22_14_port, 
      REGISTERS_22_13_port, REGISTERS_22_12_port, REGISTERS_22_11_port, 
      REGISTERS_22_10_port, REGISTERS_22_9_port, REGISTERS_22_8_port, 
      REGISTERS_22_7_port, REGISTERS_22_6_port, REGISTERS_22_5_port, 
      REGISTERS_22_4_port, REGISTERS_22_3_port, REGISTERS_22_2_port, 
      REGISTERS_22_1_port, REGISTERS_22_0_port, REGISTERS_23_31_port, 
      REGISTERS_23_30_port, REGISTERS_23_29_port, REGISTERS_23_28_port, 
      REGISTERS_23_27_port, REGISTERS_23_26_port, REGISTERS_23_25_port, 
      REGISTERS_23_24_port, REGISTERS_23_23_port, REGISTERS_23_22_port, 
      REGISTERS_23_21_port, REGISTERS_23_20_port, REGISTERS_23_19_port, 
      REGISTERS_23_18_port, REGISTERS_23_17_port, REGISTERS_23_16_port, 
      REGISTERS_23_15_port, REGISTERS_23_14_port, REGISTERS_23_13_port, 
      REGISTERS_23_12_port, REGISTERS_23_11_port, REGISTERS_23_10_port, 
      REGISTERS_23_9_port, REGISTERS_23_8_port, REGISTERS_23_7_port, 
      REGISTERS_23_6_port, REGISTERS_23_5_port, REGISTERS_23_4_port, 
      REGISTERS_23_3_port, REGISTERS_23_2_port, REGISTERS_23_1_port, 
      REGISTERS_23_0_port, REGISTERS_24_31_port, REGISTERS_24_30_port, 
      REGISTERS_24_29_port, REGISTERS_24_28_port, REGISTERS_24_27_port, 
      REGISTERS_24_26_port, REGISTERS_24_25_port, REGISTERS_24_24_port, 
      REGISTERS_24_23_port, REGISTERS_24_22_port, REGISTERS_24_21_port, 
      REGISTERS_24_20_port, REGISTERS_24_19_port, REGISTERS_24_18_port, 
      REGISTERS_24_17_port, REGISTERS_24_16_port, REGISTERS_24_15_port, 
      REGISTERS_24_14_port, REGISTERS_24_13_port, REGISTERS_24_12_port, 
      REGISTERS_24_11_port, REGISTERS_24_10_port, REGISTERS_24_9_port, 
      REGISTERS_24_8_port, REGISTERS_24_7_port, REGISTERS_24_6_port, 
      REGISTERS_24_5_port, REGISTERS_24_4_port, REGISTERS_24_3_port, 
      REGISTERS_24_2_port, REGISTERS_24_1_port, REGISTERS_24_0_port, 
      REGISTERS_25_31_port, REGISTERS_25_30_port, REGISTERS_25_29_port, 
      REGISTERS_25_28_port, REGISTERS_25_27_port, REGISTERS_25_26_port, 
      REGISTERS_25_25_port, REGISTERS_25_24_port, REGISTERS_25_23_port, 
      REGISTERS_25_22_port, REGISTERS_25_21_port, REGISTERS_25_20_port, 
      REGISTERS_25_19_port, REGISTERS_25_18_port, REGISTERS_25_17_port, 
      REGISTERS_25_16_port, REGISTERS_25_15_port, REGISTERS_25_14_port, 
      REGISTERS_25_13_port, REGISTERS_25_12_port, REGISTERS_25_11_port, 
      REGISTERS_25_10_port, REGISTERS_25_9_port, REGISTERS_25_8_port, 
      REGISTERS_25_7_port, REGISTERS_25_6_port, REGISTERS_25_5_port, 
      REGISTERS_25_4_port, REGISTERS_25_3_port, REGISTERS_25_2_port, 
      REGISTERS_25_1_port, REGISTERS_25_0_port, REGISTERS_26_31_port, 
      REGISTERS_26_30_port, REGISTERS_26_29_port, REGISTERS_26_28_port, 
      REGISTERS_26_27_port, REGISTERS_26_26_port, REGISTERS_26_25_port, 
      REGISTERS_26_24_port, REGISTERS_26_23_port, REGISTERS_26_22_port, 
      REGISTERS_26_21_port, REGISTERS_26_20_port, REGISTERS_26_19_port, 
      REGISTERS_26_18_port, REGISTERS_26_17_port, REGISTERS_26_16_port, 
      REGISTERS_26_15_port, REGISTERS_26_14_port, REGISTERS_26_13_port, 
      REGISTERS_26_12_port, REGISTERS_26_11_port, REGISTERS_26_10_port, 
      REGISTERS_26_9_port, REGISTERS_26_8_port, REGISTERS_26_7_port, 
      REGISTERS_26_6_port, REGISTERS_26_5_port, REGISTERS_26_4_port, 
      REGISTERS_26_3_port, REGISTERS_26_2_port, REGISTERS_26_1_port, 
      REGISTERS_26_0_port, REGISTERS_27_31_port, REGISTERS_27_30_port, 
      REGISTERS_27_29_port, REGISTERS_27_28_port, REGISTERS_27_27_port, 
      REGISTERS_27_26_port, REGISTERS_27_25_port, REGISTERS_27_24_port, 
      REGISTERS_27_23_port, REGISTERS_27_22_port, REGISTERS_27_21_port, 
      REGISTERS_27_20_port, REGISTERS_27_19_port, REGISTERS_27_18_port, 
      REGISTERS_27_17_port, REGISTERS_27_16_port, REGISTERS_27_15_port, 
      REGISTERS_27_14_port, REGISTERS_27_13_port, REGISTERS_27_12_port, 
      REGISTERS_27_11_port, REGISTERS_27_10_port, REGISTERS_27_9_port, 
      REGISTERS_27_8_port, REGISTERS_27_7_port, REGISTERS_27_6_port, 
      REGISTERS_27_5_port, REGISTERS_27_4_port, REGISTERS_27_3_port, 
      REGISTERS_27_2_port, REGISTERS_27_1_port, REGISTERS_27_0_port, 
      REGISTERS_28_31_port, REGISTERS_28_30_port, REGISTERS_28_29_port, 
      REGISTERS_28_28_port, REGISTERS_28_27_port, REGISTERS_28_26_port, 
      REGISTERS_28_25_port, REGISTERS_28_24_port, REGISTERS_28_23_port, 
      REGISTERS_28_22_port, REGISTERS_28_21_port, REGISTERS_28_20_port, 
      REGISTERS_28_19_port, REGISTERS_28_18_port, REGISTERS_28_17_port, 
      REGISTERS_28_16_port, REGISTERS_28_15_port, REGISTERS_28_14_port, 
      REGISTERS_28_13_port, REGISTERS_28_12_port, REGISTERS_28_11_port, 
      REGISTERS_28_10_port, REGISTERS_28_9_port, REGISTERS_28_8_port, 
      REGISTERS_28_7_port, REGISTERS_28_6_port, REGISTERS_28_5_port, 
      REGISTERS_28_4_port, REGISTERS_28_3_port, REGISTERS_28_2_port, 
      REGISTERS_28_1_port, REGISTERS_28_0_port, REGISTERS_29_31_port, 
      REGISTERS_29_30_port, REGISTERS_29_29_port, REGISTERS_29_28_port, 
      REGISTERS_29_27_port, REGISTERS_29_26_port, REGISTERS_29_25_port, 
      REGISTERS_29_24_port, REGISTERS_29_23_port, REGISTERS_29_22_port, 
      REGISTERS_29_21_port, REGISTERS_29_20_port, REGISTERS_29_19_port, 
      REGISTERS_29_18_port, REGISTERS_29_17_port, REGISTERS_29_16_port, 
      REGISTERS_29_15_port, REGISTERS_29_14_port, REGISTERS_29_13_port, 
      REGISTERS_29_12_port, REGISTERS_29_11_port, REGISTERS_29_10_port, 
      REGISTERS_29_9_port, REGISTERS_29_8_port, REGISTERS_29_7_port, 
      REGISTERS_29_6_port, REGISTERS_29_5_port, REGISTERS_29_4_port, 
      REGISTERS_29_3_port, REGISTERS_29_2_port, REGISTERS_29_1_port, 
      REGISTERS_29_0_port, REGISTERS_30_31_port, REGISTERS_30_30_port, 
      REGISTERS_30_29_port, REGISTERS_30_28_port, REGISTERS_30_27_port, 
      REGISTERS_30_26_port, REGISTERS_30_25_port, REGISTERS_30_24_port, 
      REGISTERS_30_23_port, REGISTERS_30_22_port, REGISTERS_30_21_port, 
      REGISTERS_30_20_port, REGISTERS_30_19_port, REGISTERS_30_18_port, 
      REGISTERS_30_17_port, REGISTERS_30_16_port, REGISTERS_30_15_port, 
      REGISTERS_30_14_port, REGISTERS_30_13_port, REGISTERS_30_12_port, 
      REGISTERS_30_11_port, REGISTERS_30_10_port, REGISTERS_30_9_port, 
      REGISTERS_30_8_port, REGISTERS_30_7_port, REGISTERS_30_6_port, 
      REGISTERS_30_5_port, REGISTERS_30_4_port, REGISTERS_30_3_port, 
      REGISTERS_30_2_port, REGISTERS_30_1_port, REGISTERS_30_0_port, 
      REGISTERS_31_31_port, REGISTERS_31_30_port, REGISTERS_31_29_port, 
      REGISTERS_31_28_port, REGISTERS_31_27_port, REGISTERS_31_26_port, 
      REGISTERS_31_25_port, REGISTERS_31_24_port, REGISTERS_31_23_port, 
      REGISTERS_31_22_port, REGISTERS_31_21_port, REGISTERS_31_20_port, 
      REGISTERS_31_19_port, REGISTERS_31_18_port, REGISTERS_31_17_port, 
      REGISTERS_31_16_port, REGISTERS_31_15_port, REGISTERS_31_14_port, 
      REGISTERS_31_13_port, REGISTERS_31_12_port, REGISTERS_31_11_port, 
      REGISTERS_31_10_port, REGISTERS_31_9_port, REGISTERS_31_8_port, 
      REGISTERS_31_7_port, REGISTERS_31_6_port, REGISTERS_31_5_port, 
      REGISTERS_31_4_port, REGISTERS_31_3_port, REGISTERS_31_2_port, 
      REGISTERS_31_1_port, REGISTERS_31_0_port, REGISTERS_32_31_port, 
      REGISTERS_32_30_port, REGISTERS_32_29_port, REGISTERS_32_28_port, 
      REGISTERS_32_27_port, REGISTERS_32_26_port, REGISTERS_32_25_port, 
      REGISTERS_32_24_port, REGISTERS_32_23_port, REGISTERS_32_22_port, 
      REGISTERS_32_21_port, REGISTERS_32_20_port, REGISTERS_32_19_port, 
      REGISTERS_32_18_port, REGISTERS_32_17_port, REGISTERS_32_16_port, 
      REGISTERS_32_15_port, REGISTERS_32_14_port, REGISTERS_32_13_port, 
      REGISTERS_32_12_port, REGISTERS_32_11_port, REGISTERS_32_10_port, 
      REGISTERS_32_9_port, REGISTERS_32_8_port, REGISTERS_32_7_port, 
      REGISTERS_32_6_port, REGISTERS_32_5_port, REGISTERS_32_4_port, 
      REGISTERS_32_3_port, REGISTERS_32_2_port, REGISTERS_32_1_port, 
      REGISTERS_32_0_port, REGISTERS_33_31_port, REGISTERS_33_30_port, 
      REGISTERS_33_29_port, REGISTERS_33_28_port, REGISTERS_33_27_port, 
      REGISTERS_33_26_port, REGISTERS_33_25_port, REGISTERS_33_24_port, 
      REGISTERS_33_23_port, REGISTERS_33_22_port, REGISTERS_33_21_port, 
      REGISTERS_33_20_port, REGISTERS_33_19_port, REGISTERS_33_18_port, 
      REGISTERS_33_17_port, REGISTERS_33_16_port, REGISTERS_33_15_port, 
      REGISTERS_33_14_port, REGISTERS_33_13_port, REGISTERS_33_12_port, 
      REGISTERS_33_11_port, REGISTERS_33_10_port, REGISTERS_33_9_port, 
      REGISTERS_33_8_port, REGISTERS_33_7_port, REGISTERS_33_6_port, 
      REGISTERS_33_5_port, REGISTERS_33_4_port, REGISTERS_33_3_port, 
      REGISTERS_33_2_port, REGISTERS_33_1_port, REGISTERS_33_0_port, 
      REGISTERS_34_31_port, REGISTERS_34_30_port, REGISTERS_34_29_port, 
      REGISTERS_34_28_port, REGISTERS_34_27_port, REGISTERS_34_26_port, 
      REGISTERS_34_25_port, REGISTERS_34_24_port, REGISTERS_34_23_port, 
      REGISTERS_34_22_port, REGISTERS_34_21_port, REGISTERS_34_20_port, 
      REGISTERS_34_19_port, REGISTERS_34_18_port, REGISTERS_34_17_port, 
      REGISTERS_34_16_port, REGISTERS_34_15_port, REGISTERS_34_14_port, 
      REGISTERS_34_13_port, REGISTERS_34_12_port, REGISTERS_34_11_port, 
      REGISTERS_34_10_port, REGISTERS_34_9_port, REGISTERS_34_8_port, 
      REGISTERS_34_7_port, REGISTERS_34_6_port, REGISTERS_34_5_port, 
      REGISTERS_34_4_port, REGISTERS_34_3_port, REGISTERS_34_2_port, 
      REGISTERS_34_1_port, REGISTERS_34_0_port, REGISTERS_35_31_port, 
      REGISTERS_35_30_port, REGISTERS_35_29_port, REGISTERS_35_28_port, 
      REGISTERS_35_27_port, REGISTERS_35_26_port, REGISTERS_35_25_port, 
      REGISTERS_35_24_port, REGISTERS_35_23_port, REGISTERS_35_22_port, 
      REGISTERS_35_21_port, REGISTERS_35_20_port, REGISTERS_35_19_port, 
      REGISTERS_35_18_port, REGISTERS_35_17_port, REGISTERS_35_16_port, 
      REGISTERS_35_15_port, REGISTERS_35_14_port, REGISTERS_35_13_port, 
      REGISTERS_35_12_port, REGISTERS_35_11_port, REGISTERS_35_10_port, 
      REGISTERS_35_9_port, REGISTERS_35_8_port, REGISTERS_35_7_port, 
      REGISTERS_35_6_port, REGISTERS_35_5_port, REGISTERS_35_4_port, 
      REGISTERS_35_3_port, REGISTERS_35_2_port, REGISTERS_35_1_port, 
      REGISTERS_35_0_port, REGISTERS_36_31_port, REGISTERS_36_30_port, 
      REGISTERS_36_29_port, REGISTERS_36_28_port, REGISTERS_36_27_port, 
      REGISTERS_36_26_port, REGISTERS_36_25_port, REGISTERS_36_24_port, 
      REGISTERS_36_23_port, REGISTERS_36_22_port, REGISTERS_36_21_port, 
      REGISTERS_36_20_port, REGISTERS_36_19_port, REGISTERS_36_18_port, 
      REGISTERS_36_17_port, REGISTERS_36_16_port, REGISTERS_36_15_port, 
      REGISTERS_36_14_port, REGISTERS_36_13_port, REGISTERS_36_12_port, 
      REGISTERS_36_11_port, REGISTERS_36_10_port, REGISTERS_36_9_port, 
      REGISTERS_36_8_port, REGISTERS_36_7_port, REGISTERS_36_6_port, 
      REGISTERS_36_5_port, REGISTERS_36_4_port, REGISTERS_36_3_port, 
      REGISTERS_36_2_port, REGISTERS_36_1_port, REGISTERS_36_0_port, 
      REGISTERS_37_31_port, REGISTERS_37_30_port, REGISTERS_37_29_port, 
      REGISTERS_37_28_port, REGISTERS_37_27_port, REGISTERS_37_26_port, 
      REGISTERS_37_25_port, REGISTERS_37_24_port, REGISTERS_37_23_port, 
      REGISTERS_37_22_port, REGISTERS_37_21_port, REGISTERS_37_20_port, 
      REGISTERS_37_19_port, REGISTERS_37_18_port, REGISTERS_37_17_port, 
      REGISTERS_37_16_port, REGISTERS_37_15_port, REGISTERS_37_14_port, 
      REGISTERS_37_13_port, REGISTERS_37_12_port, REGISTERS_37_11_port, 
      REGISTERS_37_10_port, REGISTERS_37_9_port, REGISTERS_37_8_port, 
      REGISTERS_37_7_port, REGISTERS_37_6_port, REGISTERS_37_5_port, 
      REGISTERS_37_4_port, REGISTERS_37_3_port, REGISTERS_37_2_port, 
      REGISTERS_37_1_port, REGISTERS_37_0_port, REGISTERS_38_31_port, 
      REGISTERS_38_30_port, REGISTERS_38_29_port, REGISTERS_38_28_port, 
      REGISTERS_38_27_port, REGISTERS_38_26_port, REGISTERS_38_25_port, 
      REGISTERS_38_24_port, REGISTERS_38_23_port, REGISTERS_38_22_port, 
      REGISTERS_38_21_port, REGISTERS_38_20_port, REGISTERS_38_19_port, 
      REGISTERS_38_18_port, REGISTERS_38_17_port, REGISTERS_38_16_port, 
      REGISTERS_38_15_port, REGISTERS_38_14_port, REGISTERS_38_13_port, 
      REGISTERS_38_12_port, REGISTERS_38_11_port, REGISTERS_38_10_port, 
      REGISTERS_38_9_port, REGISTERS_38_8_port, REGISTERS_38_7_port, 
      REGISTERS_38_6_port, REGISTERS_38_5_port, REGISTERS_38_4_port, 
      REGISTERS_38_3_port, REGISTERS_38_2_port, REGISTERS_38_1_port, 
      REGISTERS_38_0_port, REGISTERS_39_31_port, REGISTERS_39_30_port, 
      REGISTERS_39_29_port, REGISTERS_39_28_port, REGISTERS_39_27_port, 
      REGISTERS_39_26_port, REGISTERS_39_25_port, REGISTERS_39_24_port, 
      REGISTERS_39_23_port, REGISTERS_39_22_port, REGISTERS_39_21_port, 
      REGISTERS_39_20_port, REGISTERS_39_19_port, REGISTERS_39_18_port, 
      REGISTERS_39_17_port, REGISTERS_39_16_port, REGISTERS_39_15_port, 
      REGISTERS_39_14_port, REGISTERS_39_13_port, REGISTERS_39_12_port, 
      REGISTERS_39_11_port, REGISTERS_39_10_port, REGISTERS_39_9_port, 
      REGISTERS_39_8_port, REGISTERS_39_7_port, REGISTERS_39_6_port, 
      REGISTERS_39_5_port, REGISTERS_39_4_port, REGISTERS_39_3_port, 
      REGISTERS_39_2_port, REGISTERS_39_1_port, REGISTERS_39_0_port, 
      REGISTERS_40_31_port, REGISTERS_40_30_port, REGISTERS_40_29_port, 
      REGISTERS_40_28_port, REGISTERS_40_27_port, REGISTERS_40_26_port, 
      REGISTERS_40_25_port, REGISTERS_40_24_port, REGISTERS_40_23_port, 
      REGISTERS_40_22_port, REGISTERS_40_21_port, REGISTERS_40_20_port, 
      REGISTERS_40_19_port, REGISTERS_40_18_port, REGISTERS_40_17_port, 
      REGISTERS_40_16_port, REGISTERS_40_15_port, REGISTERS_40_14_port, 
      REGISTERS_40_13_port, REGISTERS_40_12_port, REGISTERS_40_11_port, 
      REGISTERS_40_10_port, REGISTERS_40_9_port, REGISTERS_40_8_port, 
      REGISTERS_40_7_port, REGISTERS_40_6_port, REGISTERS_40_5_port, 
      REGISTERS_40_4_port, REGISTERS_40_3_port, REGISTERS_40_2_port, 
      REGISTERS_40_1_port, REGISTERS_40_0_port, REGISTERS_41_31_port, 
      REGISTERS_41_30_port, REGISTERS_41_29_port, REGISTERS_41_28_port, 
      REGISTERS_41_27_port, REGISTERS_41_26_port, REGISTERS_41_25_port, 
      REGISTERS_41_24_port, REGISTERS_41_23_port, REGISTERS_41_22_port, 
      REGISTERS_41_21_port, REGISTERS_41_20_port, REGISTERS_41_19_port, 
      REGISTERS_41_18_port, REGISTERS_41_17_port, REGISTERS_41_16_port, 
      REGISTERS_41_15_port, REGISTERS_41_14_port, REGISTERS_41_13_port, 
      REGISTERS_41_12_port, REGISTERS_41_11_port, REGISTERS_41_10_port, 
      REGISTERS_41_9_port, REGISTERS_41_8_port, REGISTERS_41_7_port, 
      REGISTERS_41_6_port, REGISTERS_41_5_port, REGISTERS_41_4_port, 
      REGISTERS_41_3_port, REGISTERS_41_2_port, REGISTERS_41_1_port, 
      REGISTERS_41_0_port, REGISTERS_42_31_port, REGISTERS_42_30_port, 
      REGISTERS_42_29_port, REGISTERS_42_28_port, REGISTERS_42_27_port, 
      REGISTERS_42_26_port, REGISTERS_42_25_port, REGISTERS_42_24_port, 
      REGISTERS_42_23_port, REGISTERS_42_22_port, REGISTERS_42_21_port, 
      REGISTERS_42_20_port, REGISTERS_42_19_port, REGISTERS_42_18_port, 
      REGISTERS_42_17_port, REGISTERS_42_16_port, REGISTERS_42_15_port, 
      REGISTERS_42_14_port, REGISTERS_42_13_port, REGISTERS_42_12_port, 
      REGISTERS_42_11_port, REGISTERS_42_10_port, REGISTERS_42_9_port, 
      REGISTERS_42_8_port, REGISTERS_42_7_port, REGISTERS_42_6_port, 
      REGISTERS_42_5_port, REGISTERS_42_4_port, REGISTERS_42_3_port, 
      REGISTERS_42_2_port, REGISTERS_42_1_port, REGISTERS_42_0_port, 
      REGISTERS_43_31_port, REGISTERS_43_30_port, REGISTERS_43_29_port, 
      REGISTERS_43_28_port, REGISTERS_43_27_port, REGISTERS_43_26_port, 
      REGISTERS_43_25_port, REGISTERS_43_24_port, REGISTERS_43_23_port, 
      REGISTERS_43_22_port, REGISTERS_43_21_port, REGISTERS_43_20_port, 
      REGISTERS_43_19_port, REGISTERS_43_18_port, REGISTERS_43_17_port, 
      REGISTERS_43_16_port, REGISTERS_43_15_port, REGISTERS_43_14_port, 
      REGISTERS_43_13_port, REGISTERS_43_12_port, REGISTERS_43_11_port, 
      REGISTERS_43_10_port, REGISTERS_43_9_port, REGISTERS_43_8_port, 
      REGISTERS_43_7_port, REGISTERS_43_6_port, REGISTERS_43_5_port, 
      REGISTERS_43_4_port, REGISTERS_43_3_port, REGISTERS_43_2_port, 
      REGISTERS_43_1_port, REGISTERS_43_0_port, REGISTERS_44_31_port, 
      REGISTERS_44_30_port, REGISTERS_44_29_port, REGISTERS_44_28_port, 
      REGISTERS_44_27_port, REGISTERS_44_26_port, REGISTERS_44_25_port, 
      REGISTERS_44_24_port, REGISTERS_44_23_port, REGISTERS_44_22_port, 
      REGISTERS_44_21_port, REGISTERS_44_20_port, REGISTERS_44_19_port, 
      REGISTERS_44_18_port, REGISTERS_44_17_port, REGISTERS_44_16_port, 
      REGISTERS_44_15_port, REGISTERS_44_14_port, REGISTERS_44_13_port, 
      REGISTERS_44_12_port, REGISTERS_44_11_port, REGISTERS_44_10_port, 
      REGISTERS_44_9_port, REGISTERS_44_8_port, REGISTERS_44_7_port, 
      REGISTERS_44_6_port, REGISTERS_44_5_port, REGISTERS_44_4_port, 
      REGISTERS_44_3_port, REGISTERS_44_2_port, REGISTERS_44_1_port, 
      REGISTERS_44_0_port, REGISTERS_45_31_port, REGISTERS_45_30_port, 
      REGISTERS_45_29_port, REGISTERS_45_28_port, REGISTERS_45_27_port, 
      REGISTERS_45_26_port, REGISTERS_45_25_port, REGISTERS_45_24_port, 
      REGISTERS_45_23_port, REGISTERS_45_22_port, REGISTERS_45_21_port, 
      REGISTERS_45_20_port, REGISTERS_45_19_port, REGISTERS_45_18_port, 
      REGISTERS_45_17_port, REGISTERS_45_16_port, REGISTERS_45_15_port, 
      REGISTERS_45_14_port, REGISTERS_45_13_port, REGISTERS_45_12_port, 
      REGISTERS_45_11_port, REGISTERS_45_10_port, REGISTERS_45_9_port, 
      REGISTERS_45_8_port, REGISTERS_45_7_port, REGISTERS_45_6_port, 
      REGISTERS_45_5_port, REGISTERS_45_4_port, REGISTERS_45_3_port, 
      REGISTERS_45_2_port, REGISTERS_45_1_port, REGISTERS_45_0_port, 
      REGISTERS_46_31_port, REGISTERS_46_30_port, REGISTERS_46_29_port, 
      REGISTERS_46_28_port, REGISTERS_46_27_port, REGISTERS_46_26_port, 
      REGISTERS_46_25_port, REGISTERS_46_24_port, REGISTERS_46_23_port, 
      REGISTERS_46_22_port, REGISTERS_46_21_port, REGISTERS_46_20_port, 
      REGISTERS_46_19_port, REGISTERS_46_18_port, REGISTERS_46_17_port, 
      REGISTERS_46_16_port, REGISTERS_46_15_port, REGISTERS_46_14_port, 
      REGISTERS_46_13_port, REGISTERS_46_12_port, REGISTERS_46_11_port, 
      REGISTERS_46_10_port, REGISTERS_46_9_port, REGISTERS_46_8_port, 
      REGISTERS_46_7_port, REGISTERS_46_6_port, REGISTERS_46_5_port, 
      REGISTERS_46_4_port, REGISTERS_46_3_port, REGISTERS_46_2_port, 
      REGISTERS_46_1_port, REGISTERS_46_0_port, REGISTERS_47_31_port, 
      REGISTERS_47_30_port, REGISTERS_47_29_port, REGISTERS_47_28_port, 
      REGISTERS_47_27_port, REGISTERS_47_26_port, REGISTERS_47_25_port, 
      REGISTERS_47_24_port, REGISTERS_47_23_port, REGISTERS_47_22_port, 
      REGISTERS_47_21_port, REGISTERS_47_20_port, REGISTERS_47_19_port, 
      REGISTERS_47_18_port, REGISTERS_47_17_port, REGISTERS_47_16_port, 
      REGISTERS_47_15_port, REGISTERS_47_14_port, REGISTERS_47_13_port, 
      REGISTERS_47_12_port, REGISTERS_47_11_port, REGISTERS_47_10_port, 
      REGISTERS_47_9_port, REGISTERS_47_8_port, REGISTERS_47_7_port, 
      REGISTERS_47_6_port, REGISTERS_47_5_port, REGISTERS_47_4_port, 
      REGISTERS_47_3_port, REGISTERS_47_2_port, REGISTERS_47_1_port, 
      REGISTERS_47_0_port, REGISTERS_48_31_port, REGISTERS_48_30_port, 
      REGISTERS_48_29_port, REGISTERS_48_28_port, REGISTERS_48_27_port, 
      REGISTERS_48_26_port, REGISTERS_48_25_port, REGISTERS_48_24_port, 
      REGISTERS_48_23_port, REGISTERS_48_22_port, REGISTERS_48_21_port, 
      REGISTERS_48_20_port, REGISTERS_48_19_port, REGISTERS_48_18_port, 
      REGISTERS_48_17_port, REGISTERS_48_16_port, REGISTERS_48_15_port, 
      REGISTERS_48_14_port, REGISTERS_48_13_port, REGISTERS_48_12_port, 
      REGISTERS_48_11_port, REGISTERS_48_10_port, REGISTERS_48_9_port, 
      REGISTERS_48_8_port, REGISTERS_48_7_port, REGISTERS_48_6_port, 
      REGISTERS_48_5_port, REGISTERS_48_4_port, REGISTERS_48_3_port, 
      REGISTERS_48_2_port, REGISTERS_48_1_port, REGISTERS_48_0_port, 
      REGISTERS_49_31_port, REGISTERS_49_30_port, REGISTERS_49_29_port, 
      REGISTERS_49_28_port, REGISTERS_49_27_port, REGISTERS_49_26_port, 
      REGISTERS_49_25_port, REGISTERS_49_24_port, REGISTERS_49_23_port, 
      REGISTERS_49_22_port, REGISTERS_49_21_port, REGISTERS_49_20_port, 
      REGISTERS_49_19_port, REGISTERS_49_18_port, REGISTERS_49_17_port, 
      REGISTERS_49_16_port, REGISTERS_49_15_port, REGISTERS_49_14_port, 
      REGISTERS_49_13_port, REGISTERS_49_12_port, REGISTERS_49_11_port, 
      REGISTERS_49_10_port, REGISTERS_49_9_port, REGISTERS_49_8_port, 
      REGISTERS_49_7_port, REGISTERS_49_6_port, REGISTERS_49_5_port, 
      REGISTERS_49_4_port, REGISTERS_49_3_port, REGISTERS_49_2_port, 
      REGISTERS_49_1_port, REGISTERS_49_0_port, REGISTERS_50_31_port, 
      REGISTERS_50_30_port, REGISTERS_50_29_port, REGISTERS_50_28_port, 
      REGISTERS_50_27_port, REGISTERS_50_26_port, REGISTERS_50_25_port, 
      REGISTERS_50_24_port, REGISTERS_50_23_port, REGISTERS_50_22_port, 
      REGISTERS_50_21_port, REGISTERS_50_20_port, REGISTERS_50_19_port, 
      REGISTERS_50_18_port, REGISTERS_50_17_port, REGISTERS_50_16_port, 
      REGISTERS_50_15_port, REGISTERS_50_14_port, REGISTERS_50_13_port, 
      REGISTERS_50_12_port, REGISTERS_50_11_port, REGISTERS_50_10_port, 
      REGISTERS_50_9_port, REGISTERS_50_8_port, REGISTERS_50_7_port, 
      REGISTERS_50_6_port, REGISTERS_50_5_port, REGISTERS_50_4_port, 
      REGISTERS_50_3_port, REGISTERS_50_2_port, REGISTERS_50_1_port, 
      REGISTERS_50_0_port, REGISTERS_51_31_port, REGISTERS_51_30_port, 
      REGISTERS_51_29_port, REGISTERS_51_28_port, REGISTERS_51_27_port, 
      REGISTERS_51_26_port, REGISTERS_51_25_port, REGISTERS_51_24_port, 
      REGISTERS_51_23_port, REGISTERS_51_22_port, REGISTERS_51_21_port, 
      REGISTERS_51_20_port, REGISTERS_51_19_port, REGISTERS_51_18_port, 
      REGISTERS_51_17_port, REGISTERS_51_16_port, REGISTERS_51_15_port, 
      REGISTERS_51_14_port, REGISTERS_51_13_port, REGISTERS_51_12_port, 
      REGISTERS_51_11_port, REGISTERS_51_10_port, REGISTERS_51_9_port, 
      REGISTERS_51_8_port, REGISTERS_51_7_port, REGISTERS_51_6_port, 
      REGISTERS_51_5_port, REGISTERS_51_4_port, REGISTERS_51_3_port, 
      REGISTERS_51_2_port, REGISTERS_51_1_port, REGISTERS_51_0_port, 
      REGISTERS_52_31_port, REGISTERS_52_30_port, REGISTERS_52_29_port, 
      REGISTERS_52_28_port, REGISTERS_52_27_port, REGISTERS_52_26_port, 
      REGISTERS_52_25_port, REGISTERS_52_24_port, REGISTERS_52_23_port, 
      REGISTERS_52_22_port, REGISTERS_52_21_port, REGISTERS_52_20_port, 
      REGISTERS_52_19_port, REGISTERS_52_18_port, REGISTERS_52_17_port, 
      REGISTERS_52_16_port, REGISTERS_52_15_port, REGISTERS_52_14_port, 
      REGISTERS_52_13_port, REGISTERS_52_12_port, REGISTERS_52_11_port, 
      REGISTERS_52_10_port, REGISTERS_52_9_port, REGISTERS_52_8_port, 
      REGISTERS_52_7_port, REGISTERS_52_6_port, REGISTERS_52_5_port, 
      REGISTERS_52_4_port, REGISTERS_52_3_port, REGISTERS_52_2_port, 
      REGISTERS_52_1_port, REGISTERS_52_0_port, REGISTERS_53_31_port, 
      REGISTERS_53_30_port, REGISTERS_53_29_port, REGISTERS_53_28_port, 
      REGISTERS_53_27_port, REGISTERS_53_26_port, REGISTERS_53_25_port, 
      REGISTERS_53_24_port, REGISTERS_53_23_port, REGISTERS_53_22_port, 
      REGISTERS_53_21_port, REGISTERS_53_20_port, REGISTERS_53_19_port, 
      REGISTERS_53_18_port, REGISTERS_53_17_port, REGISTERS_53_16_port, 
      REGISTERS_53_15_port, REGISTERS_53_14_port, REGISTERS_53_13_port, 
      REGISTERS_53_12_port, REGISTERS_53_11_port, REGISTERS_53_10_port, 
      REGISTERS_53_9_port, REGISTERS_53_8_port, REGISTERS_53_7_port, 
      REGISTERS_53_6_port, REGISTERS_53_5_port, REGISTERS_53_4_port, 
      REGISTERS_53_3_port, REGISTERS_53_2_port, REGISTERS_53_1_port, 
      REGISTERS_53_0_port, REGISTERS_54_31_port, REGISTERS_54_30_port, 
      REGISTERS_54_29_port, REGISTERS_54_28_port, REGISTERS_54_27_port, 
      REGISTERS_54_26_port, REGISTERS_54_25_port, REGISTERS_54_24_port, 
      REGISTERS_54_23_port, REGISTERS_54_22_port, REGISTERS_54_21_port, 
      REGISTERS_54_20_port, REGISTERS_54_19_port, REGISTERS_54_18_port, 
      REGISTERS_54_17_port, REGISTERS_54_16_port, REGISTERS_54_15_port, 
      REGISTERS_54_14_port, REGISTERS_54_13_port, REGISTERS_54_12_port, 
      REGISTERS_54_11_port, REGISTERS_54_10_port, REGISTERS_54_9_port, 
      REGISTERS_54_8_port, REGISTERS_54_7_port, REGISTERS_54_6_port, 
      REGISTERS_54_5_port, REGISTERS_54_4_port, REGISTERS_54_3_port, 
      REGISTERS_54_2_port, REGISTERS_54_1_port, REGISTERS_54_0_port, 
      REGISTERS_55_31_port, REGISTERS_55_30_port, REGISTERS_55_29_port, 
      REGISTERS_55_28_port, REGISTERS_55_27_port, REGISTERS_55_26_port, 
      REGISTERS_55_25_port, REGISTERS_55_24_port, REGISTERS_55_23_port, 
      REGISTERS_55_22_port, REGISTERS_55_21_port, REGISTERS_55_20_port, 
      REGISTERS_55_19_port, REGISTERS_55_18_port, REGISTERS_55_17_port, 
      REGISTERS_55_16_port, REGISTERS_55_15_port, REGISTERS_55_14_port, 
      REGISTERS_55_13_port, REGISTERS_55_12_port, REGISTERS_55_11_port, 
      REGISTERS_55_10_port, REGISTERS_55_9_port, REGISTERS_55_8_port, 
      REGISTERS_55_7_port, REGISTERS_55_6_port, REGISTERS_55_5_port, 
      REGISTERS_55_4_port, REGISTERS_55_3_port, REGISTERS_55_2_port, 
      REGISTERS_55_1_port, REGISTERS_55_0_port, REGISTERS_56_31_port, 
      REGISTERS_56_30_port, REGISTERS_56_29_port, REGISTERS_56_28_port, 
      REGISTERS_56_27_port, REGISTERS_56_26_port, REGISTERS_56_25_port, 
      REGISTERS_56_24_port, REGISTERS_56_23_port, REGISTERS_56_22_port, 
      REGISTERS_56_21_port, REGISTERS_56_20_port, REGISTERS_56_19_port, 
      REGISTERS_56_18_port, REGISTERS_56_17_port, REGISTERS_56_16_port, 
      REGISTERS_56_15_port, REGISTERS_56_14_port, REGISTERS_56_13_port, 
      REGISTERS_56_12_port, REGISTERS_56_11_port, REGISTERS_56_10_port, 
      REGISTERS_56_9_port, REGISTERS_56_8_port, REGISTERS_56_7_port, 
      REGISTERS_56_6_port, REGISTERS_56_5_port, REGISTERS_56_4_port, 
      REGISTERS_56_3_port, REGISTERS_56_2_port, REGISTERS_56_1_port, 
      REGISTERS_56_0_port, REGISTERS_57_31_port, REGISTERS_57_30_port, 
      REGISTERS_57_29_port, REGISTERS_57_28_port, REGISTERS_57_27_port, 
      REGISTERS_57_26_port, REGISTERS_57_25_port, REGISTERS_57_24_port, 
      REGISTERS_57_23_port, REGISTERS_57_22_port, REGISTERS_57_21_port, 
      REGISTERS_57_20_port, REGISTERS_57_19_port, REGISTERS_57_18_port, 
      REGISTERS_57_17_port, REGISTERS_57_16_port, REGISTERS_57_15_port, 
      REGISTERS_57_14_port, REGISTERS_57_13_port, REGISTERS_57_12_port, 
      REGISTERS_57_11_port, REGISTERS_57_10_port, REGISTERS_57_9_port, 
      REGISTERS_57_8_port, REGISTERS_57_7_port, REGISTERS_57_6_port, 
      REGISTERS_57_5_port, REGISTERS_57_4_port, REGISTERS_57_3_port, 
      REGISTERS_57_2_port, REGISTERS_57_1_port, REGISTERS_57_0_port, 
      REGISTERS_58_31_port, REGISTERS_58_30_port, REGISTERS_58_29_port, 
      REGISTERS_58_28_port, REGISTERS_58_27_port, REGISTERS_58_26_port, 
      REGISTERS_58_25_port, REGISTERS_58_24_port, REGISTERS_58_23_port, 
      REGISTERS_58_22_port, REGISTERS_58_21_port, REGISTERS_58_20_port, 
      REGISTERS_58_19_port, REGISTERS_58_18_port, REGISTERS_58_17_port, 
      REGISTERS_58_16_port, REGISTERS_58_15_port, REGISTERS_58_14_port, 
      REGISTERS_58_13_port, REGISTERS_58_12_port, REGISTERS_58_11_port, 
      REGISTERS_58_10_port, REGISTERS_58_9_port, REGISTERS_58_8_port, 
      REGISTERS_58_7_port, REGISTERS_58_6_port, REGISTERS_58_5_port, 
      REGISTERS_58_4_port, REGISTERS_58_3_port, REGISTERS_58_2_port, 
      REGISTERS_58_1_port, REGISTERS_58_0_port, REGISTERS_59_31_port, 
      REGISTERS_59_30_port, REGISTERS_59_29_port, REGISTERS_59_28_port, 
      REGISTERS_59_27_port, REGISTERS_59_26_port, REGISTERS_59_25_port, 
      REGISTERS_59_24_port, REGISTERS_59_23_port, REGISTERS_59_22_port, 
      REGISTERS_59_21_port, REGISTERS_59_20_port, REGISTERS_59_19_port, 
      REGISTERS_59_18_port, REGISTERS_59_17_port, REGISTERS_59_16_port, 
      REGISTERS_59_15_port, REGISTERS_59_14_port, REGISTERS_59_13_port, 
      REGISTERS_59_12_port, REGISTERS_59_11_port, REGISTERS_59_10_port, 
      REGISTERS_59_9_port, REGISTERS_59_8_port, REGISTERS_59_7_port, 
      REGISTERS_59_6_port, REGISTERS_59_5_port, REGISTERS_59_4_port, 
      REGISTERS_59_3_port, REGISTERS_59_2_port, REGISTERS_59_1_port, 
      REGISTERS_59_0_port, REGISTERS_60_31_port, REGISTERS_60_30_port, 
      REGISTERS_60_29_port, REGISTERS_60_28_port, REGISTERS_60_27_port, 
      REGISTERS_60_26_port, REGISTERS_60_25_port, REGISTERS_60_24_port, 
      REGISTERS_60_23_port, REGISTERS_60_22_port, REGISTERS_60_21_port, 
      REGISTERS_60_20_port, REGISTERS_60_19_port, REGISTERS_60_18_port, 
      REGISTERS_60_17_port, REGISTERS_60_16_port, REGISTERS_60_15_port, 
      REGISTERS_60_14_port, REGISTERS_60_13_port, REGISTERS_60_12_port, 
      REGISTERS_60_11_port, REGISTERS_60_10_port, REGISTERS_60_9_port, 
      REGISTERS_60_8_port, REGISTERS_60_7_port, REGISTERS_60_6_port, 
      REGISTERS_60_5_port, REGISTERS_60_4_port, REGISTERS_60_3_port, 
      REGISTERS_60_2_port, REGISTERS_60_1_port, REGISTERS_60_0_port, 
      REGISTERS_61_31_port, REGISTERS_61_30_port, REGISTERS_61_29_port, 
      REGISTERS_61_28_port, REGISTERS_61_27_port, REGISTERS_61_26_port, 
      REGISTERS_61_25_port, REGISTERS_61_24_port, REGISTERS_61_23_port, 
      REGISTERS_61_22_port, REGISTERS_61_21_port, REGISTERS_61_20_port, 
      REGISTERS_61_19_port, REGISTERS_61_18_port, REGISTERS_61_17_port, 
      REGISTERS_61_16_port, REGISTERS_61_15_port, REGISTERS_61_14_port, 
      REGISTERS_61_13_port, REGISTERS_61_12_port, REGISTERS_61_11_port, 
      REGISTERS_61_10_port, REGISTERS_61_9_port, REGISTERS_61_8_port, 
      REGISTERS_61_7_port, REGISTERS_61_6_port, REGISTERS_61_5_port, 
      REGISTERS_61_4_port, REGISTERS_61_3_port, REGISTERS_61_2_port, 
      REGISTERS_61_1_port, REGISTERS_61_0_port, REGISTERS_62_31_port, 
      REGISTERS_62_30_port, REGISTERS_62_29_port, REGISTERS_62_28_port, 
      REGISTERS_62_27_port, REGISTERS_62_26_port, REGISTERS_62_25_port, 
      REGISTERS_62_24_port, REGISTERS_62_23_port, REGISTERS_62_22_port, 
      REGISTERS_62_21_port, REGISTERS_62_20_port, REGISTERS_62_19_port, 
      REGISTERS_62_18_port, REGISTERS_62_17_port, REGISTERS_62_16_port, 
      REGISTERS_62_15_port, REGISTERS_62_14_port, REGISTERS_62_13_port, 
      REGISTERS_62_12_port, REGISTERS_62_11_port, REGISTERS_62_10_port, 
      REGISTERS_62_9_port, REGISTERS_62_8_port, REGISTERS_62_7_port, 
      REGISTERS_62_6_port, REGISTERS_62_5_port, REGISTERS_62_4_port, 
      REGISTERS_62_3_port, REGISTERS_62_2_port, REGISTERS_62_1_port, 
      REGISTERS_62_0_port, REGISTERS_63_31_port, REGISTERS_63_30_port, 
      REGISTERS_63_29_port, REGISTERS_63_28_port, REGISTERS_63_27_port, 
      REGISTERS_63_26_port, REGISTERS_63_25_port, REGISTERS_63_24_port, 
      REGISTERS_63_23_port, REGISTERS_63_22_port, REGISTERS_63_21_port, 
      REGISTERS_63_20_port, REGISTERS_63_19_port, REGISTERS_63_18_port, 
      REGISTERS_63_17_port, REGISTERS_63_16_port, REGISTERS_63_15_port, 
      REGISTERS_63_14_port, REGISTERS_63_13_port, REGISTERS_63_12_port, 
      REGISTERS_63_11_port, REGISTERS_63_10_port, REGISTERS_63_9_port, 
      REGISTERS_63_8_port, REGISTERS_63_7_port, REGISTERS_63_6_port, 
      REGISTERS_63_5_port, REGISTERS_63_4_port, REGISTERS_63_3_port, 
      REGISTERS_63_2_port, REGISTERS_63_1_port, REGISTERS_63_0_port, N17, N18, 
      N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33
      , N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, 
      N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62
      , N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, 
      N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91
      , N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103, N104, 
      N105, N106, N107, N108, N109, N110, N111, N112, N113, N114, N115, N116, 
      N117, N118, N119, N120, N121, N122, N123, N124, N125, N126, N127, N128, 
      N129, N130, N131, N132, N133, N134, N135, N136, N137, N138, N139, N140, 
      N141, N142, N143, N144, N145, N146, N147, N148, N149, N150, N151, N152, 
      N153, N154, N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, 
      N165, N166, N167, N168, N169, N170, N171, N172, N173, N174, N175, N176, 
      N177, N178, N179, N180, N181, N182, N183, N184, N185, N186, N187, N188, 
      N189, N190, N191, N192, N193, N194, N195, N196, N197, N198, N199, N200, 
      N201, N202, N203, N204, N205, N206, N207, N208, N209, N210, N211, N212, 
      N213, N214, N215, N216, N217, N218, N219, N220, N221, N222, N223, N224, 
      N225, N226, N227, N228, N229, N230, N231, N232, N233, N234, N235, N236, 
      N237, N238, N239, N240, N241, N242, N243, N244, N245, N246, N247, N248, 
      N249, N250, N251, N252, N253, N254, N255, N256, N257, N258, N259, N260, 
      N261, N262, N263, N264, N265, N266, N267, N268, N269, N270, N271, N272, 
      N273, N274, N275, N276, N277, N278, N279, N280, N281, N282, N283, N284, 
      N285, N286, N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, 
      N297, N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308, 
      N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319, N320, 
      N321, N322, N323, N324, N325, N326, N327, N328, N329, N330, N331, N332, 
      N333, N334, N335, N336, N337, N338, N339, N340, N341, N342, N343, N344, 
      N345, N346, N347, N348, N349, N350, N351, N352, N353, N354, N355, N356, 
      N357, N358, N359, N360, N361, N362, N363, N364, N365, N366, N367, N368, 
      N369, N370, N371, N372, N373, N374, N375, N376, N377, N378, N379, N380, 
      N381, N382, N383, N384, N385, N386, N387, N388, N389, N390, N391, N392, 
      N393, N394, N395, N396, N397, N398, N399, N400, N401, N402, N403, N404, 
      N405, N406, N407, N408, N409, N410, N411, N412, N413, N414, N415, N416, 
      N417, N418, N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, 
      N429, N430, N431, N432, N433, N434, N435, N436, N437, N438, N439, N440, 
      N441, N442, N443, N444, N445, N446, N447, N448, N449, N450, N451, N452, 
      N453, N454, N455, N456, N457, N458, N459, N460, N461, N462, N463, N464, 
      N465, N466, N467, N468, N469, N470, N471, N472, N473, N474, N475, N476, 
      N477, N478, N479, N480, N481, N482, N483, N484, N485, N486, N487, N488, 
      N489, N490, N491, N492, N493, N494, N495, N496, N497, N498, N499, N500, 
      N501, N502, N503, N504, N505, N506, N507, N508, N509, N510, N511, N512, 
      N513, N514, N515, N516, N517, N518, N519, N520, N521, N522, N523, N524, 
      N525, N526, N527, N528, N529, N530, N531, N532, N533, N534, N535, N536, 
      N537, N538, N539, N540, N541, N542, N543, N544, N545, N546, N547, N548, 
      N549, N550, N551, N552, N553, N554, N555, N556, N557, N558, N559, N560, 
      N561, N562, N563, N564, N565, N566, N567, N568, N569, N570, N571, N572, 
      N573, N574, N575, N576, N577, N578, N579, N580, N581, N582, N583, N584, 
      N585, N586, N587, N588, N589, N590, N591, N592, N593, N594, N595, N596, 
      N597, N598, N599, N600, N601, N602, N603, N604, N605, N606, N607, N608, 
      N609, N610, N611, N612, N613, N614, N615, N616, N617, N618, N619, N620, 
      N621, N622, N623, N624, N625, N626, N627, N628, N629, N630, N631, N632, 
      N633, N634, N635, N636, N637, N638, N639, N640, N641, N642, N643, N644, 
      N645, N646, N647, N648, N649, N650, N651, N652, N653, N654, N655, N656, 
      N657, N658, N659, N660, N661, N662, N663, N664, N665, N666, N667, N668, 
      N669, N670, N671, N672, N673, N674, N675, N676, N677, N678, N679, N680, 
      N681, N682, N683, N684, N685, N686, N687, N688, N689, N690, N691, N692, 
      N693, N694, N695, N696, N697, N698, N699, N700, N701, N702, N703, N704, 
      N705, N706, N707, N708, N709, N710, N711, N712, N713, N714, N715, N716, 
      N717, N718, N719, N720, N721, N722, N723, N724, N725, N726, N727, N728, 
      N729, n_1000, n_1001, n_1002, n_1003, n_1004, n_1005, n_1006, n_1007, 
      n_1008, n_1009, n_1010, n_1011, n_1012, n_1013, n_1014, n_1015, n_1016, 
      n_1017, n_1018, n_1019, n_1020, n_1021, n_1022, n_1023, n_1024, n_1025, 
      n_1026, n_1027, n_1028, n_1029, n_1030, n_1031, n_1032, n_1033, n_1034, 
      n_1035, n_1036, n_1037, n_1038, n_1039, n_1040, n_1041, n_1042, n_1043, 
      n_1044, n_1045, n_1046, n_1047, n_1048, n_1049, n_1050, n_1051, n_1052, 
      n_1053, n_1054, n_1055, n_1056, n_1057, n_1058, n_1059, n_1060, n_1061, 
      n_1062, n_1063, n_1064, n_1065, n_1066, n_1067, n_1068, n_1069, n_1070, 
      n_1071, n_1072, n_1073, n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, 
      n_1080, n_1081, n_1082, n_1083, n_1084, n_1085, n_1086, n_1087, n_1088, 
      n_1089, n_1090, n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, 
      n_1098, n_1099, n_1100, n_1101, n_1102, n_1103, n_1104, n_1105, n_1106, 
      n_1107, n_1108, n_1109, n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, 
      n_1116, n_1117, n_1118, n_1119, n_1120, n_1121, n_1122, n_1123, n_1124, 
      n_1125, n_1126, n_1127, n_1128, n_1129, n_1130, n_1131, n_1132, n_1133, 
      n_1134, n_1135, n_1136, n_1137, n_1138, n_1139, n_1140, n_1141, n_1142, 
      n_1143, n_1144, n_1145, n_1146, n_1147, n_1148, n_1149, n_1150, n_1151, 
      n_1152, n_1153, n_1154, n_1155, n_1156, n_1157, n_1158, n_1159, n_1160, 
      n_1161, n_1162, n_1163, n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, 
      n_1170, n_1171, n_1172, n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, 
      n_1179, n_1180, n_1181, n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, 
      n_1188, n_1189, n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, n_1196, 
      n_1197, n_1198, n_1199, n_1200, n_1201, n_1202, n_1203, n_1204, n_1205, 
      n_1206, n_1207, n_1208, n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, 
      n_1215, n_1216, n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, 
      n_1224, n_1225, n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, n_1232, 
      n_1233, n_1234, n_1235, n_1236, n_1237, n_1238, n_1239, n_1240, n_1241, 
      n_1242, n_1243, n_1244, n_1245, n_1246, n_1247, n_1248, n_1249, n_1250, 
      n_1251, n_1252, n_1253, n_1254, n_1255, n_1256, n_1257, n_1258, n_1259, 
      n_1260, n_1261, n_1262, n_1263, n_1264, n_1265, n_1266, n_1267, n_1268, 
      n_1269, n_1270, n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, 
      n_1278, n_1279, n_1280, n_1281, n_1282, n_1283, n_1284, n_1285, n_1286, 
      n_1287, n_1288, n_1289, n_1290, n_1291, n_1292, n_1293, n_1294, n_1295, 
      n_1296, n_1297, n_1298, n_1299, n_1300, n_1301, n_1302, n_1303, n_1304, 
      n_1305, n_1306, n_1307, n_1308, n_1309, n_1310, n_1311, n_1312, n_1313, 
      n_1314, n_1315, n_1316, n_1317, n_1318, n_1319, n_1320, n_1321, n_1322, 
      n_1323, n_1324, n_1325, n_1326, n_1327, n_1328, n_1329, n_1330, n_1331, 
      n_1332, n_1333, n_1334, n_1335, n_1336, n_1337, n_1338, n_1339, n_1340, 
      n_1341, n_1342, n_1343, n_1344, n_1345, n_1346, n_1347, n_1348, n_1349, 
      n_1350, n_1351, n_1352, n_1353, n_1354, n_1355, n_1356, n_1357, n_1358, 
      n_1359, n_1360, n_1361, n_1362, n_1363, n_1364, n_1365, n_1366, n_1367, 
      n_1368, n_1369, n_1370, n_1371, n_1372, n_1373, n_1374, n_1375, n_1376, 
      n_1377, n_1378, n_1379, n_1380, n_1381, n_1382, n_1383, n_1384, n_1385, 
      n_1386, n_1387, n_1388, n_1389, n_1390, n_1391, n_1392, n_1393, n_1394, 
      n_1395, n_1396, n_1397, n_1398, n_1399, n_1400, n_1401, n_1402, n_1403, 
      n_1404, n_1405, n_1406, n_1407, n_1408, n_1409, n_1410, n_1411, n_1412, 
      n_1413, n_1414, n_1415, n_1416, n_1417, n_1418, n_1419, n_1420, n_1421, 
      n_1422, n_1423, n_1424, n_1425, n_1426, n_1427, n_1428, n_1429, n_1430, 
      n_1431, n_1432, n_1433, n_1434, n_1435, n_1436, n_1437, n_1438, n_1439, 
      n_1440, n_1441, n_1442, n_1443, n_1444, n_1445, n_1446, n_1447, n_1448, 
      n_1449, n_1450, n_1451, n_1452, n_1453, n_1454, n_1455, n_1456, n_1457, 
      n_1458, n_1459, n_1460, n_1461, n_1462, n_1463, n_1464, n_1465, n_1466, 
      n_1467, n_1468, n_1469, n_1470, n_1471, n_1472, n_1473, n_1474, n_1475, 
      n_1476, n_1477, n_1478, n_1479, n_1480, n_1481, n_1482, n_1483, n_1484, 
      n_1485, n_1486, n_1487, n_1488, n_1489, n_1490, n_1491, n_1492, n_1493, 
      n_1494, n_1495, n_1496, n_1497, n_1498, n_1499, n_1500, n_1501, n_1502, 
      n_1503, n_1504, n_1505, n_1506, n_1507, n_1508, n_1509, n_1510, n_1511, 
      n_1512, n_1513, n_1514, n_1515, n_1516, n_1517, n_1518, n_1519, n_1520, 
      n_1521, n_1522, n_1523, n_1524, n_1525, n_1526, n_1527, n_1528, n_1529, 
      n_1530, n_1531, n_1532, n_1533, n_1534, n_1535, n_1536, n_1537, n_1538, 
      n_1539, n_1540, n_1541, n_1542, n_1543, n_1544, n_1545, n_1546, n_1547, 
      n_1548, n_1549, n_1550, n_1551, n_1552, n_1553, n_1554, n_1555, n_1556, 
      n_1557, n_1558, n_1559, n_1560, n_1561, n_1562, n_1563, n_1564, n_1565, 
      n_1566, n_1567, n_1568, n_1569, n_1570, n_1571, n_1572, n_1573, n_1574, 
      n_1575, n_1576, n_1577, n_1578, n_1579, n_1580, n_1581, n_1582, n_1583, 
      n_1584, n_1585, n_1586, n_1587, n_1588, n_1589, n_1590, n_1591, n_1592, 
      n_1593, n_1594, n_1595, n_1596, n_1597, n_1598, n_1599, n_1600, n_1601, 
      n_1602, n_1603, n_1604, n_1605, n_1606, n_1607, n_1608, n_1609, n_1610, 
      n_1611, n_1612, n_1613, n_1614, n_1615, n_1616, n_1617, n_1618, n_1619, 
      n_1620, n_1621, n_1622, n_1623, n_1624, n_1625, n_1626, n_1627, n_1628, 
      n_1629, n_1630, n_1631, n_1632, n_1633, n_1634, n_1635, n_1636, n_1637, 
      n_1638, n_1639, n_1640, n_1641, n_1642, n_1643, n_1644, n_1645, n_1646, 
      n_1647, n_1648, n_1649, n_1650, n_1651, n_1652, n_1653, n_1654, n_1655, 
      n_1656, n_1657, n_1658, n_1659, n_1660, n_1661, n_1662, n_1663, n_1664, 
      n_1665, n_1666, n_1667, n_1668, n_1669, n_1670, n_1671, n_1672, n_1673, 
      n_1674, n_1675, n_1676, n_1677, n_1678, n_1679, n_1680, n_1681, n_1682, 
      n_1683, n_1684, n_1685, n_1686, n_1687, n_1688, n_1689, n_1690, n_1691, 
      n_1692, n_1693, n_1694, n_1695, n_1696, n_1697, n_1698, n_1699, n_1700, 
      n_1701, n_1702, n_1703, n_1704, n_1705, n_1706, n_1707, n_1708, n_1709, 
      n_1710, n_1711, n_1712, n_1713, n_1714, n_1715, n_1716, n_1717, n_1718, 
      n_1719, n_1720, n_1721, n_1722, n_1723, n_1724, n_1725, n_1726, n_1727, 
      n_1728, n_1729, n_1730, n_1731, n_1732, n_1733, n_1734, n_1735, n_1736, 
      n_1737, n_1738, n_1739, n_1740, n_1741, n_1742, n_1743, n_1744, n_1745, 
      n_1746, n_1747, n_1748, n_1749, n_1750, n_1751, n_1752, n_1753, n_1754, 
      n_1755, n_1756, n_1757, n_1758, n_1759, n_1760, n_1761, n_1762, n_1763, 
      n_1764, n_1765, n_1766, n_1767, n_1768, n_1769, n_1770, n_1771, n_1772, 
      n_1773, n_1774, n_1775, n_1776, n_1777, n_1778, n_1779, n_1780, n_1781, 
      n_1782, n_1783, n_1784, n_1785, n_1786, n_1787, n_1788, n_1789, n_1790, 
      n_1791, n_1792, n_1793, n_1794, n_1795, n_1796, n_1797, n_1798, n_1799, 
      n_1800, n_1801, n_1802, n_1803, n_1804, n_1805, n_1806, n_1807, n_1808, 
      n_1809, n_1810, n_1811, n_1812, n_1813, n_1814, n_1815, n_1816, n_1817, 
      n_1818, n_1819, n_1820, n_1821, n_1822, n_1823, n_1824, n_1825, n_1826, 
      n_1827, n_1828, n_1829, n_1830, n_1831, n_1832, n_1833, n_1834, n_1835, 
      n_1836, n_1837, n_1838, n_1839, n_1840, n_1841, n_1842, n_1843, n_1844, 
      n_1845, n_1846, n_1847, n_1848, n_1849, n_1850, n_1851, n_1852, n_1853, 
      n_1854, n_1855, n_1856, n_1857, n_1858, n_1859, n_1860, n_1861, n_1862, 
      n_1863, n_1864, n_1865, n_1866, n_1867, n_1868, n_1869, n_1870, n_1871, 
      n_1872, n_1873, n_1874, n_1875, n_1876, n_1877, n_1878, n_1879, n_1880, 
      n_1881, n_1882, n_1883, n_1884, n_1885, n_1886, n_1887, n_1888, n_1889, 
      n_1890, n_1891, n_1892, n_1893, n_1894, n_1895, n_1896, n_1897, n_1898, 
      n_1899, n_1900, n_1901, n_1902, n_1903, n_1904, n_1905, n_1906, n_1907, 
      n_1908, n_1909, n_1910, n_1911, n_1912, n_1913, n_1914, n_1915, n_1916, 
      n_1917, n_1918, n_1919, n_1920, n_1921, n_1922, n_1923, n_1924, n_1925, 
      n_1926, n_1927, n_1928, n_1929, n_1930, n_1931, n_1932, n_1933, n_1934, 
      n_1935, n_1936, n_1937, n_1938, n_1939, n_1940, n_1941, n_1942, n_1943, 
      n_1944, n_1945, n_1946, n_1947, n_1948, n_1949, n_1950, n_1951, n_1952, 
      n_1953, n_1954, n_1955, n_1956, n_1957, n_1958, n_1959, n_1960, n_1961, 
      n_1962, n_1963, n_1964, n_1965, n_1966, n_1967, n_1968, n_1969, n_1970, 
      n_1971, n_1972, n_1973, n_1974, n_1975, n_1976, n_1977, n_1978, n_1979, 
      n_1980, n_1981, n_1982, n_1983, n_1984, n_1985, n_1986, n_1987, n_1988, 
      n_1989, n_1990, n_1991, n_1992, n_1993, n_1994, n_1995, n_1996, n_1997, 
      n_1998, n_1999, n_2000, n_2001, n_2002, n_2003, n_2004, n_2005, n_2006, 
      n_2007, n_2008, n_2009, n_2010, n_2011, n_2012, n_2013, n_2014, n_2015, 
      n_2016, n_2017, n_2018, n_2019, n_2020, n_2021, n_2022, n_2023, n_2024, 
      n_2025, n_2026, n_2027, n_2028, n_2029, n_2030, n_2031, n_2032, n_2033, 
      n_2034, n_2035, n_2036, n_2037, n_2038, n_2039, n_2040, n_2041, n_2042, 
      n_2043, n_2044, n_2045, n_2046, n_2047, n_2048, n_2049, n_2050, n_2051, 
      n_2052, n_2053, n_2054, n_2055, n_2056, n_2057, n_2058, n_2059, n_2060, 
      n_2061, n_2062, n_2063, n_2064, n_2065, n_2066, n_2067, n_2068, n_2069, 
      n_2070, n_2071, n_2072, n_2073, n_2074, n_2075, n_2076, n_2077, n_2078, 
      n_2079, n_2080, n_2081, n_2082, n_2083, n_2084, n_2085, n_2086, n_2087, 
      n_2088, n_2089, n_2090, n_2091, n_2092, n_2093, n_2094, n_2095, n_2096, 
      n_2097, n_2098, n_2099, n_2100, n_2101, n_2102, n_2103, n_2104, n_2105, 
      n_2106, n_2107, n_2108, n_2109, n_2110, n_2111, n_2112, n_2113, n_2114, 
      n_2115, n_2116, n_2117, n_2118, n_2119, n_2120, n_2121, n_2122, n_2123, 
      n_2124, n_2125, n_2126, n_2127, n_2128, n_2129, n_2130, n_2131, n_2132, 
      n_2133, n_2134, n_2135, n_2136, n_2137, n_2138, n_2139, n_2140, n_2141, 
      n_2142, n_2143, n_2144, n_2145, n_2146, n_2147, n_2148, n_2149, n_2150, 
      n_2151, n_2152, n_2153, n_2154, n_2155, n_2156, n_2157, n_2158, n_2159, 
      n_2160, n_2161, n_2162, n_2163, n_2164, n_2165, n_2166, n_2167, n_2168, 
      n_2169, n_2170, n_2171, n_2172, n_2173, n_2174, n_2175, n_2176, n_2177, 
      n_2178, n_2179, n_2180, n_2181, n_2182, n_2183, n_2184, n_2185, n_2186, 
      n_2187, n_2188, n_2189, n_2190, n_2191, n_2192, n_2193, n_2194, n_2195, 
      n_2196, n_2197, n_2198, n_2199, n_2200, n_2201, n_2202, n_2203, n_2204, 
      n_2205, n_2206, n_2207, n_2208, n_2209, n_2210, n_2211, n_2212, n_2213, 
      n_2214, n_2215, n_2216, n_2217, n_2218, n_2219, n_2220, n_2221, n_2222, 
      n_2223, n_2224, n_2225, n_2226, n_2227, n_2228, n_2229, n_2230, n_2231, 
      n_2232, n_2233, n_2234, n_2235, n_2236, n_2237, n_2238, n_2239, n_2240, 
      n_2241, n_2242, n_2243, n_2244, n_2245, n_2246, n_2247, n_2248, n_2249, 
      n_2250, n_2251, n_2252, n_2253, n_2254, n_2255, n_2256, n_2257, n_2258, 
      n_2259, n_2260, n_2261, n_2262, n_2263, n_2264, n_2265, n_2266, n_2267, 
      n_2268, n_2269, n_2270, n_2271, n_2272, n_2273, n_2274, n_2275, n_2276, 
      n_2277, n_2278, n_2279, n_2280, n_2281, n_2282, n_2283, n_2284, n_2285, 
      n_2286, n_2287, n_2288, n_2289, n_2290, n_2291, n_2292, n_2293, n_2294, 
      n_2295, n_2296, n_2297, n_2298, n_2299, n_2300, n_2301, n_2302, n_2303, 
      n_2304, n_2305, n_2306, n_2307, n_2308, n_2309, n_2310, n_2311, n_2312, 
      n_2313, n_2314, n_2315, n_2316, n_2317, n_2318, n_2319, n_2320, n_2321, 
      n_2322, n_2323, n_2324, n_2325, n_2326, n_2327, n_2328, n_2329, n_2330, 
      n_2331, n_2332, n_2333, n_2334, n_2335, n_2336, n_2337, n_2338, n_2339, 
      n_2340, n_2341, n_2342, n_2343, n_2344, n_2345, n_2346, n_2347, n_2348, 
      n_2349, n_2350, n_2351, n_2352, n_2353, n_2354, n_2355, n_2356, n_2357, 
      n_2358, n_2359, n_2360, n_2361, n_2362, n_2363, n_2364, n_2365, n_2366, 
      n_2367, n_2368, n_2369, n_2370, n_2371, n_2372, n_2373, n_2374, n_2375, 
      n_2376, n_2377, n_2378, n_2379, n_2380, n_2381, n_2382, n_2383, n_2384, 
      n_2385, n_2386, n_2387, n_2388, n_2389, n_2390, n_2391, n_2392, n_2393, 
      n_2394, n_2395, n_2396, n_2397, n_2398, n_2399, n_2400, n_2401, n_2402, 
      n_2403, n_2404, n_2405, n_2406, n_2407, n_2408, n_2409, n_2410, n_2411, 
      n_2412, n_2413, n_2414, n_2415, n_2416, n_2417, n_2418, n_2419, n_2420, 
      n_2421, n_2422, n_2423, n_2424, n_2425, n_2426, n_2427, n_2428, n_2429, 
      n_2430, n_2431, n_2432, n_2433, n_2434, n_2435, n_2436, n_2437, n_2438, 
      n_2439, n_2440, n_2441, n_2442, n_2443, n_2444, n_2445, n_2446, n_2447, 
      n_2448, n_2449, n_2450, n_2451, n_2452, n_2453, n_2454, n_2455, n_2456, 
      n_2457, n_2458, n_2459, n_2460, n_2461, n_2462, n_2463, n_2464, n_2465, 
      n_2466, n_2467, n_2468, n_2469, n_2470, n_2471, n_2472, n_2473, n_2474, 
      n_2475, n_2476, n_2477, n_2478, n_2479, n_2480, n_2481, n_2482, n_2483, 
      n_2484, n_2485, n_2486, n_2487, n_2488, n_2489, n_2490, n_2491, n_2492, 
      n_2493, n_2494, n_2495, n_2496, n_2497, n_2498, n_2499, n_2500, n_2501, 
      n_2502, n_2503, n_2504, n_2505, n_2506, n_2507, n_2508, n_2509, n_2510, 
      n_2511, n_2512, n_2513, n_2514, n_2515, n_2516, n_2517, n_2518, n_2519, 
      n_2520, n_2521, n_2522, n_2523, n_2524, n_2525, n_2526, n_2527, n_2528, 
      n_2529, n_2530, n_2531, n_2532, n_2533, n_2534, n_2535, n_2536, n_2537, 
      n_2538, n_2539, n_2540, n_2541, n_2542, n_2543, n_2544, n_2545, n_2546, 
      n_2547, n_2548, n_2549, n_2550, n_2551, n_2552, n_2553, n_2554, n_2555, 
      n_2556, n_2557, n_2558, n_2559, n_2560, n_2561, n_2562, n_2563, n_2564, 
      n_2565, n_2566, n_2567, n_2568, n_2569, n_2570, n_2571, n_2572, n_2573, 
      n_2574, n_2575, n_2576, n_2577, n_2578, n_2579, n_2580, n_2581, n_2582, 
      n_2583, n_2584, n_2585, n_2586, n_2587, n_2588, n_2589, n_2590, n_2591, 
      n_2592, n_2593, n_2594, n_2595, n_2596, n_2597, n_2598, n_2599, n_2600, 
      n_2601, n_2602, n_2603, n_2604, n_2605, n_2606, n_2607, n_2608, n_2609, 
      n_2610, n_2611, n_2612, n_2613, n_2614, n_2615, n_2616, n_2617, n_2618, 
      n_2619, n_2620, n_2621, n_2622, n_2623, n_2624, n_2625, n_2626, n_2627, 
      n_2628, n_2629, n_2630, n_2631, n_2632, n_2633, n_2634, n_2635, n_2636, 
      n_2637, n_2638, n_2639, n_2640, n_2641, n_2642, n_2643, n_2644, n_2645, 
      n_2646, n_2647, n_2648, n_2649, n_2650, n_2651, n_2652, n_2653, n_2654, 
      n_2655, n_2656, n_2657, n_2658, n_2659, n_2660, n_2661, n_2662, n_2663, 
      n_2664, n_2665, n_2666, n_2667, n_2668, n_2669, n_2670, n_2671, n_2672, 
      n_2673, n_2674, n_2675, n_2676, n_2677, n_2678, n_2679, n_2680, n_2681, 
      n_2682, n_2683, n_2684, n_2685, n_2686, n_2687, n_2688, n_2689, n_2690, 
      n_2691, n_2692, n_2693, n_2694, n_2695, n_2696, n_2697, n_2698, n_2699, 
      n_2700, n_2701, n_2702, n_2703, n_2704, n_2705, n_2706, n_2707, n_2708, 
      n_2709, n_2710, n_2711, n_2712, n_2713, n_2714, n_2715, n_2716, n_2717, 
      n_2718, n_2719, n_2720, n_2721, n_2722, n_2723, n_2724, n_2725, n_2726, 
      n_2727, n_2728, n_2729, n_2730, n_2731, n_2732, n_2733, n_2734, n_2735, 
      n_2736, n_2737, n_2738, n_2739, n_2740, n_2741, n_2742, n_2743, n_2744, 
      n_2745, n_2746, n_2747, n_2748, n_2749, n_2750, n_2751, n_2752, n_2753, 
      n_2754, n_2755, n_2756, n_2757, n_2758, n_2759, n_2760, n_2761, n_2762, 
      n_2763, n_2764, n_2765, n_2766, n_2767, n_2768, n_2769, n_2770, n_2771, 
      n_2772, n_2773, n_2774, n_2775, n_2776, n_2777, n_2778, n_2779, n_2780, 
      n_2781, n_2782, n_2783, n_2784, n_2785, n_2786, n_2787, n_2788, n_2789, 
      n_2790, n_2791, n_2792, n_2793, n_2794, n_2795, n_2796, n_2797, n_2798, 
      n_2799, n_2800, n_2801, n_2802, n_2803, n_2804, n_2805, n_2806, n_2807, 
      n_2808, n_2809, n_2810, n_2811, n_2812, n_2813, n_2814, n_2815, n_2816, 
      n_2817, n_2818, n_2819, n_2820, n_2821, n_2822, n_2823, n_2824, n_2825, 
      n_2826, n_2827, n_2828, n_2829, n_2830, n_2831, n_2832, n_2833, n_2834, 
      n_2835, n_2836, n_2837, n_2838, n_2839, n_2840, n_2841, n_2842, n_2843, 
      n_2844, n_2845, n_2846, n_2847, n_2848, n_2849, n_2850, n_2851, n_2852, 
      n_2853, n_2854, n_2855, n_2856, n_2857, n_2858, n_2859, n_2860, n_2861, 
      n_2862, n_2863, n_2864, n_2865, n_2866, n_2867, n_2868, n_2869, n_2870, 
      n_2871, n_2872, n_2873, n_2874, n_2875, n_2876, n_2877, n_2878, n_2879, 
      n_2880, n_2881, n_2882, n_2883, n_2884, n_2885, n_2886, n_2887, n_2888, 
      n_2889, n_2890, n_2891, n_2892, n_2893, n_2894, n_2895, n_2896, n_2897, 
      n_2898, n_2899, n_2900, n_2901, n_2902, n_2903, n_2904, n_2905, n_2906, 
      n_2907, n_2908, n_2909, n_2910, n_2911, n_2912, n_2913, n_2914, n_2915, 
      n_2916, n_2917, n_2918, n_2919, n_2920, n_2921, n_2922, n_2923, n_2924, 
      n_2925, n_2926, n_2927, n_2928, n_2929, n_2930, n_2931, n_2932, n_2933, 
      n_2934, n_2935, n_2936, n_2937, n_2938, n_2939, n_2940, n_2941, n_2942, 
      n_2943, n_2944, n_2945, n_2946, n_2947, n_2948, n_2949, n_2950, n_2951, 
      n_2952, n_2953, n_2954, n_2955, n_2956, n_2957, n_2958, n_2959, n_2960, 
      n_2961, n_2962, n_2963, n_2964, n_2965, n_2966, n_2967, n_2968, n_2969, 
      n_2970, n_2971, n_2972, n_2973, n_2974, n_2975, n_2976, n_2977, n_2978, 
      n_2979, n_2980, n_2981, n_2982, n_2983, n_2984, n_2985, n_2986, n_2987, 
      n_2988, n_2989, n_2990, n_2991, n_2992, n_2993, n_2994, n_2995, n_2996, 
      n_2997, n_2998, n_2999, n_3000, n_3001, n_3002, n_3003, n_3004, n_3005, 
      n_3006, n_3007, n_3008, n_3009, n_3010, n_3011, n_3012, n_3013, n_3014, 
      n_3015, n_3016, n_3017, n_3018, n_3019, n_3020, n_3021, n_3022, n_3023, 
      n_3024, n_3025, n_3026, n_3027, n_3028, n_3029, n_3030, n_3031, n_3032, 
      n_3033, n_3034, n_3035, n_3036, n_3037, n_3038, n_3039, n_3040, n_3041, 
      n_3042, n_3043, n_3044, n_3045, n_3046, n_3047, n_3048, n_3049, n_3050, 
      n_3051, n_3052, n_3053, n_3054, n_3055, n_3056, n_3057, n_3058, n_3059, 
      n_3060, n_3061, n_3062, n_3063, n_3064, n_3065, n_3066, n_3067, n_3068, 
      n_3069, n_3070, n_3071, n_3072, n_3073, n_3074, n_3075, n_3076, n_3077, 
      n_3078, n_3079, n_3080, n_3081, n_3082, n_3083, n_3084, n_3085, n_3086, 
      n_3087, n_3088, n_3089, n_3090, n_3091, n_3092, n_3093, n_3094, n_3095, 
      n_3096, n_3097, n_3098, n_3099, n_3100, n_3101, n_3102, n_3103, n_3104, 
      n_3105, n_3106, n_3107, n_3108, n_3109, n_3110, n_3111 : std_logic;

begin
   CLK_port <= CLK;
   RD1_port <= RD1;
   RD2_port <= RD2;
   ( DATAIN_31_port, DATAIN_30_port, DATAIN_29_port, DATAIN_28_port, 
      DATAIN_27_port, DATAIN_26_port, DATAIN_25_port, DATAIN_24_port, 
      DATAIN_23_port, DATAIN_22_port, DATAIN_21_port, DATAIN_20_port, 
      DATAIN_19_port, DATAIN_18_port, DATAIN_17_port, DATAIN_16_port, 
      DATAIN_15_port, DATAIN_14_port, DATAIN_13_port, DATAIN_12_port, 
      DATAIN_11_port, DATAIN_10_port, DATAIN_9_port, DATAIN_8_port, 
      DATAIN_7_port, DATAIN_6_port, DATAIN_5_port, DATAIN_4_port, DATAIN_3_port
      , DATAIN_2_port, DATAIN_1_port, DATAIN_0_port ) <= DATAIN;
   OUT1 <= ( OUT1_31_port, OUT1_30_port, OUT1_29_port, OUT1_28_port, 
      OUT1_27_port, OUT1_26_port, OUT1_25_port, OUT1_24_port, OUT1_23_port, 
      OUT1_22_port, OUT1_21_port, OUT1_20_port, OUT1_19_port, OUT1_18_port, 
      OUT1_17_port, OUT1_16_port, OUT1_15_port, OUT1_14_port, OUT1_13_port, 
      OUT1_12_port, OUT1_11_port, OUT1_10_port, OUT1_9_port, OUT1_8_port, 
      OUT1_7_port, OUT1_6_port, OUT1_5_port, OUT1_4_port, OUT1_3_port, 
      OUT1_2_port, OUT1_1_port, OUT1_0_port );
   OUT2 <= ( OUT2_31_port, OUT2_30_port, OUT2_29_port, OUT2_28_port, 
      OUT2_27_port, OUT2_26_port, OUT2_25_port, OUT2_24_port, OUT2_23_port, 
      OUT2_22_port, OUT2_21_port, OUT2_20_port, OUT2_19_port, OUT2_18_port, 
      OUT2_17_port, OUT2_16_port, OUT2_15_port, OUT2_14_port, OUT2_13_port, 
      OUT2_12_port, OUT2_11_port, OUT2_10_port, OUT2_9_port, OUT2_8_port, 
      OUT2_7_port, OUT2_6_port, OUT2_5_port, OUT2_4_port, OUT2_3_port, 
      OUT2_2_port, OUT2_1_port, OUT2_0_port );
   
   REGISTERS_reg_0_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N178, next_state => N115, 
               clocked_on => CLK_port, Q => REGISTERS_0_31_port, QN => n_1000);
   REGISTERS_reg_0_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N178, next_state => N114, 
               clocked_on => CLK_port, Q => REGISTERS_0_30_port, QN => n_1001);
   REGISTERS_reg_0_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N178, next_state => N113, 
               clocked_on => CLK_port, Q => REGISTERS_0_29_port, QN => n_1002);
   REGISTERS_reg_0_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N178, next_state => N112, 
               clocked_on => CLK_port, Q => REGISTERS_0_28_port, QN => n_1003);
   REGISTERS_reg_0_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N178, next_state => N111, 
               clocked_on => CLK_port, Q => REGISTERS_0_27_port, QN => n_1004);
   REGISTERS_reg_0_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N178, next_state => N110, 
               clocked_on => CLK_port, Q => REGISTERS_0_26_port, QN => n_1005);
   REGISTERS_reg_0_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N178, next_state => N109, 
               clocked_on => CLK_port, Q => REGISTERS_0_25_port, QN => n_1006);
   REGISTERS_reg_0_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N178, next_state => N108, 
               clocked_on => CLK_port, Q => REGISTERS_0_24_port, QN => n_1007);
   REGISTERS_reg_0_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N178, next_state => N107, 
               clocked_on => CLK_port, Q => REGISTERS_0_23_port, QN => n_1008);
   REGISTERS_reg_0_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N178, next_state => N106, 
               clocked_on => CLK_port, Q => REGISTERS_0_22_port, QN => n_1009);
   REGISTERS_reg_0_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N178, next_state => N105, 
               clocked_on => CLK_port, Q => REGISTERS_0_21_port, QN => n_1010);
   REGISTERS_reg_0_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N178, next_state => N104, 
               clocked_on => CLK_port, Q => REGISTERS_0_20_port, QN => n_1011);
   REGISTERS_reg_0_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N178, next_state => N103, 
               clocked_on => CLK_port, Q => REGISTERS_0_19_port, QN => n_1012);
   REGISTERS_reg_0_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N178, next_state => N102, 
               clocked_on => CLK_port, Q => REGISTERS_0_18_port, QN => n_1013);
   REGISTERS_reg_0_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N178, next_state => N101, 
               clocked_on => CLK_port, Q => REGISTERS_0_17_port, QN => n_1014);
   REGISTERS_reg_0_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N178, next_state => N100, 
               clocked_on => CLK_port, Q => REGISTERS_0_16_port, QN => n_1015);
   REGISTERS_reg_0_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N178, next_state => N99, 
               clocked_on => CLK_port, Q => REGISTERS_0_15_port, QN => n_1016);
   REGISTERS_reg_0_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N178, next_state => N98, 
               clocked_on => CLK_port, Q => REGISTERS_0_14_port, QN => n_1017);
   REGISTERS_reg_0_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N178, next_state => N97, 
               clocked_on => CLK_port, Q => REGISTERS_0_13_port, QN => n_1018);
   REGISTERS_reg_0_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N178, next_state => N96, 
               clocked_on => CLK_port, Q => REGISTERS_0_12_port, QN => n_1019);
   REGISTERS_reg_0_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N178, next_state => N95, 
               clocked_on => CLK_port, Q => REGISTERS_0_11_port, QN => n_1020);
   REGISTERS_reg_0_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N178, next_state => N94, 
               clocked_on => CLK_port, Q => REGISTERS_0_10_port, QN => n_1021);
   REGISTERS_reg_0_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N178, next_state => N93, 
               clocked_on => CLK_port, Q => REGISTERS_0_9_port, QN => n_1022);
   REGISTERS_reg_0_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N178, next_state => N92, 
               clocked_on => CLK_port, Q => REGISTERS_0_8_port, QN => n_1023);
   REGISTERS_reg_0_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N178, next_state => N91, 
               clocked_on => CLK_port, Q => REGISTERS_0_7_port, QN => n_1024);
   REGISTERS_reg_0_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N178, next_state => N90, 
               clocked_on => CLK_port, Q => REGISTERS_0_6_port, QN => n_1025);
   REGISTERS_reg_0_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N178, next_state => N89, 
               clocked_on => CLK_port, Q => REGISTERS_0_5_port, QN => n_1026);
   REGISTERS_reg_0_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N178, next_state => N88, 
               clocked_on => CLK_port, Q => REGISTERS_0_4_port, QN => n_1027);
   REGISTERS_reg_0_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N178, next_state => N87, 
               clocked_on => CLK_port, Q => REGISTERS_0_3_port, QN => n_1028);
   REGISTERS_reg_0_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N178, next_state => N86, 
               clocked_on => CLK_port, Q => REGISTERS_0_2_port, QN => n_1029);
   REGISTERS_reg_0_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N178, next_state => N85, 
               clocked_on => CLK_port, Q => REGISTERS_0_1_port, QN => n_1030);
   REGISTERS_reg_0_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N178, next_state => N84, 
               clocked_on => CLK_port, Q => REGISTERS_0_0_port, QN => n_1031);
   REGISTERS_reg_1_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N177, next_state => N115, 
               clocked_on => CLK_port, Q => REGISTERS_1_31_port, QN => n_1032);
   REGISTERS_reg_1_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N177, next_state => N114, 
               clocked_on => CLK_port, Q => REGISTERS_1_30_port, QN => n_1033);
   REGISTERS_reg_1_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N177, next_state => N113, 
               clocked_on => CLK_port, Q => REGISTERS_1_29_port, QN => n_1034);
   REGISTERS_reg_1_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N177, next_state => N112, 
               clocked_on => CLK_port, Q => REGISTERS_1_28_port, QN => n_1035);
   REGISTERS_reg_1_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N177, next_state => N111, 
               clocked_on => CLK_port, Q => REGISTERS_1_27_port, QN => n_1036);
   REGISTERS_reg_1_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N177, next_state => N110, 
               clocked_on => CLK_port, Q => REGISTERS_1_26_port, QN => n_1037);
   REGISTERS_reg_1_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N177, next_state => N109, 
               clocked_on => CLK_port, Q => REGISTERS_1_25_port, QN => n_1038);
   REGISTERS_reg_1_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N177, next_state => N108, 
               clocked_on => CLK_port, Q => REGISTERS_1_24_port, QN => n_1039);
   REGISTERS_reg_1_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N177, next_state => N107, 
               clocked_on => CLK_port, Q => REGISTERS_1_23_port, QN => n_1040);
   REGISTERS_reg_1_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N177, next_state => N106, 
               clocked_on => CLK_port, Q => REGISTERS_1_22_port, QN => n_1041);
   REGISTERS_reg_1_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N177, next_state => N105, 
               clocked_on => CLK_port, Q => REGISTERS_1_21_port, QN => n_1042);
   REGISTERS_reg_1_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N177, next_state => N104, 
               clocked_on => CLK_port, Q => REGISTERS_1_20_port, QN => n_1043);
   REGISTERS_reg_1_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N177, next_state => N103, 
               clocked_on => CLK_port, Q => REGISTERS_1_19_port, QN => n_1044);
   REGISTERS_reg_1_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N177, next_state => N102, 
               clocked_on => CLK_port, Q => REGISTERS_1_18_port, QN => n_1045);
   REGISTERS_reg_1_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N177, next_state => N101, 
               clocked_on => CLK_port, Q => REGISTERS_1_17_port, QN => n_1046);
   REGISTERS_reg_1_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N177, next_state => N100, 
               clocked_on => CLK_port, Q => REGISTERS_1_16_port, QN => n_1047);
   REGISTERS_reg_1_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N177, next_state => N99, 
               clocked_on => CLK_port, Q => REGISTERS_1_15_port, QN => n_1048);
   REGISTERS_reg_1_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N177, next_state => N98, 
               clocked_on => CLK_port, Q => REGISTERS_1_14_port, QN => n_1049);
   REGISTERS_reg_1_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N177, next_state => N97, 
               clocked_on => CLK_port, Q => REGISTERS_1_13_port, QN => n_1050);
   REGISTERS_reg_1_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N177, next_state => N96, 
               clocked_on => CLK_port, Q => REGISTERS_1_12_port, QN => n_1051);
   REGISTERS_reg_1_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N177, next_state => N95, 
               clocked_on => CLK_port, Q => REGISTERS_1_11_port, QN => n_1052);
   REGISTERS_reg_1_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N177, next_state => N94, 
               clocked_on => CLK_port, Q => REGISTERS_1_10_port, QN => n_1053);
   REGISTERS_reg_1_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N177, next_state => N93, 
               clocked_on => CLK_port, Q => REGISTERS_1_9_port, QN => n_1054);
   REGISTERS_reg_1_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N177, next_state => N92, 
               clocked_on => CLK_port, Q => REGISTERS_1_8_port, QN => n_1055);
   REGISTERS_reg_1_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N177, next_state => N91, 
               clocked_on => CLK_port, Q => REGISTERS_1_7_port, QN => n_1056);
   REGISTERS_reg_1_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N177, next_state => N90, 
               clocked_on => CLK_port, Q => REGISTERS_1_6_port, QN => n_1057);
   REGISTERS_reg_1_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N177, next_state => N89, 
               clocked_on => CLK_port, Q => REGISTERS_1_5_port, QN => n_1058);
   REGISTERS_reg_1_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N177, next_state => N88, 
               clocked_on => CLK_port, Q => REGISTERS_1_4_port, QN => n_1059);
   REGISTERS_reg_1_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N177, next_state => N87, 
               clocked_on => CLK_port, Q => REGISTERS_1_3_port, QN => n_1060);
   REGISTERS_reg_1_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N177, next_state => N86, 
               clocked_on => CLK_port, Q => REGISTERS_1_2_port, QN => n_1061);
   REGISTERS_reg_1_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N177, next_state => N85, 
               clocked_on => CLK_port, Q => REGISTERS_1_1_port, QN => n_1062);
   REGISTERS_reg_1_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N177, next_state => N84, 
               clocked_on => CLK_port, Q => REGISTERS_1_0_port, QN => n_1063);
   REGISTERS_reg_2_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N176, next_state => N115, 
               clocked_on => CLK_port, Q => REGISTERS_2_31_port, QN => n_1064);
   REGISTERS_reg_2_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N176, next_state => N114, 
               clocked_on => CLK_port, Q => REGISTERS_2_30_port, QN => n_1065);
   REGISTERS_reg_2_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N176, next_state => N113, 
               clocked_on => CLK_port, Q => REGISTERS_2_29_port, QN => n_1066);
   REGISTERS_reg_2_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N176, next_state => N112, 
               clocked_on => CLK_port, Q => REGISTERS_2_28_port, QN => n_1067);
   REGISTERS_reg_2_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N176, next_state => N111, 
               clocked_on => CLK_port, Q => REGISTERS_2_27_port, QN => n_1068);
   REGISTERS_reg_2_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N176, next_state => N110, 
               clocked_on => CLK_port, Q => REGISTERS_2_26_port, QN => n_1069);
   REGISTERS_reg_2_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N176, next_state => N109, 
               clocked_on => CLK_port, Q => REGISTERS_2_25_port, QN => n_1070);
   REGISTERS_reg_2_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N176, next_state => N108, 
               clocked_on => CLK_port, Q => REGISTERS_2_24_port, QN => n_1071);
   REGISTERS_reg_2_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N176, next_state => N107, 
               clocked_on => CLK_port, Q => REGISTERS_2_23_port, QN => n_1072);
   REGISTERS_reg_2_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N176, next_state => N106, 
               clocked_on => CLK_port, Q => REGISTERS_2_22_port, QN => n_1073);
   REGISTERS_reg_2_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N176, next_state => N105, 
               clocked_on => CLK_port, Q => REGISTERS_2_21_port, QN => n_1074);
   REGISTERS_reg_2_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N176, next_state => N104, 
               clocked_on => CLK_port, Q => REGISTERS_2_20_port, QN => n_1075);
   REGISTERS_reg_2_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N176, next_state => N103, 
               clocked_on => CLK_port, Q => REGISTERS_2_19_port, QN => n_1076);
   REGISTERS_reg_2_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N176, next_state => N102, 
               clocked_on => CLK_port, Q => REGISTERS_2_18_port, QN => n_1077);
   REGISTERS_reg_2_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N176, next_state => N101, 
               clocked_on => CLK_port, Q => REGISTERS_2_17_port, QN => n_1078);
   REGISTERS_reg_2_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N176, next_state => N100, 
               clocked_on => CLK_port, Q => REGISTERS_2_16_port, QN => n_1079);
   REGISTERS_reg_2_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N176, next_state => N99, 
               clocked_on => CLK_port, Q => REGISTERS_2_15_port, QN => n_1080);
   REGISTERS_reg_2_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N176, next_state => N98, 
               clocked_on => CLK_port, Q => REGISTERS_2_14_port, QN => n_1081);
   REGISTERS_reg_2_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N176, next_state => N97, 
               clocked_on => CLK_port, Q => REGISTERS_2_13_port, QN => n_1082);
   REGISTERS_reg_2_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N176, next_state => N96, 
               clocked_on => CLK_port, Q => REGISTERS_2_12_port, QN => n_1083);
   REGISTERS_reg_2_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N176, next_state => N95, 
               clocked_on => CLK_port, Q => REGISTERS_2_11_port, QN => n_1084);
   REGISTERS_reg_2_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N176, next_state => N94, 
               clocked_on => CLK_port, Q => REGISTERS_2_10_port, QN => n_1085);
   REGISTERS_reg_2_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N176, next_state => N93, 
               clocked_on => CLK_port, Q => REGISTERS_2_9_port, QN => n_1086);
   REGISTERS_reg_2_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N176, next_state => N92, 
               clocked_on => CLK_port, Q => REGISTERS_2_8_port, QN => n_1087);
   REGISTERS_reg_2_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N176, next_state => N91, 
               clocked_on => CLK_port, Q => REGISTERS_2_7_port, QN => n_1088);
   REGISTERS_reg_2_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N176, next_state => N90, 
               clocked_on => CLK_port, Q => REGISTERS_2_6_port, QN => n_1089);
   REGISTERS_reg_2_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N176, next_state => N89, 
               clocked_on => CLK_port, Q => REGISTERS_2_5_port, QN => n_1090);
   REGISTERS_reg_2_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N176, next_state => N88, 
               clocked_on => CLK_port, Q => REGISTERS_2_4_port, QN => n_1091);
   REGISTERS_reg_2_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N176, next_state => N87, 
               clocked_on => CLK_port, Q => REGISTERS_2_3_port, QN => n_1092);
   REGISTERS_reg_2_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N176, next_state => N86, 
               clocked_on => CLK_port, Q => REGISTERS_2_2_port, QN => n_1093);
   REGISTERS_reg_2_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N176, next_state => N85, 
               clocked_on => CLK_port, Q => REGISTERS_2_1_port, QN => n_1094);
   REGISTERS_reg_2_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N176, next_state => N84, 
               clocked_on => CLK_port, Q => REGISTERS_2_0_port, QN => n_1095);
   REGISTERS_reg_3_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N175, next_state => N115, 
               clocked_on => CLK_port, Q => REGISTERS_3_31_port, QN => n_1096);
   REGISTERS_reg_3_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N175, next_state => N114, 
               clocked_on => CLK_port, Q => REGISTERS_3_30_port, QN => n_1097);
   REGISTERS_reg_3_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N175, next_state => N113, 
               clocked_on => CLK_port, Q => REGISTERS_3_29_port, QN => n_1098);
   REGISTERS_reg_3_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N175, next_state => N112, 
               clocked_on => CLK_port, Q => REGISTERS_3_28_port, QN => n_1099);
   REGISTERS_reg_3_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N175, next_state => N111, 
               clocked_on => CLK_port, Q => REGISTERS_3_27_port, QN => n_1100);
   REGISTERS_reg_3_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N175, next_state => N110, 
               clocked_on => CLK_port, Q => REGISTERS_3_26_port, QN => n_1101);
   REGISTERS_reg_3_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N175, next_state => N109, 
               clocked_on => CLK_port, Q => REGISTERS_3_25_port, QN => n_1102);
   REGISTERS_reg_3_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N175, next_state => N108, 
               clocked_on => CLK_port, Q => REGISTERS_3_24_port, QN => n_1103);
   REGISTERS_reg_3_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N175, next_state => N107, 
               clocked_on => CLK_port, Q => REGISTERS_3_23_port, QN => n_1104);
   REGISTERS_reg_3_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N175, next_state => N106, 
               clocked_on => CLK_port, Q => REGISTERS_3_22_port, QN => n_1105);
   REGISTERS_reg_3_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N175, next_state => N105, 
               clocked_on => CLK_port, Q => REGISTERS_3_21_port, QN => n_1106);
   REGISTERS_reg_3_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N175, next_state => N104, 
               clocked_on => CLK_port, Q => REGISTERS_3_20_port, QN => n_1107);
   REGISTERS_reg_3_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N175, next_state => N103, 
               clocked_on => CLK_port, Q => REGISTERS_3_19_port, QN => n_1108);
   REGISTERS_reg_3_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N175, next_state => N102, 
               clocked_on => CLK_port, Q => REGISTERS_3_18_port, QN => n_1109);
   REGISTERS_reg_3_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N175, next_state => N101, 
               clocked_on => CLK_port, Q => REGISTERS_3_17_port, QN => n_1110);
   REGISTERS_reg_3_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N175, next_state => N100, 
               clocked_on => CLK_port, Q => REGISTERS_3_16_port, QN => n_1111);
   REGISTERS_reg_3_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N175, next_state => N99, 
               clocked_on => CLK_port, Q => REGISTERS_3_15_port, QN => n_1112);
   REGISTERS_reg_3_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N175, next_state => N98, 
               clocked_on => CLK_port, Q => REGISTERS_3_14_port, QN => n_1113);
   REGISTERS_reg_3_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N175, next_state => N97, 
               clocked_on => CLK_port, Q => REGISTERS_3_13_port, QN => n_1114);
   REGISTERS_reg_3_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N175, next_state => N96, 
               clocked_on => CLK_port, Q => REGISTERS_3_12_port, QN => n_1115);
   REGISTERS_reg_3_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N175, next_state => N95, 
               clocked_on => CLK_port, Q => REGISTERS_3_11_port, QN => n_1116);
   REGISTERS_reg_3_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N175, next_state => N94, 
               clocked_on => CLK_port, Q => REGISTERS_3_10_port, QN => n_1117);
   REGISTERS_reg_3_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N175, next_state => N93, 
               clocked_on => CLK_port, Q => REGISTERS_3_9_port, QN => n_1118);
   REGISTERS_reg_3_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N175, next_state => N92, 
               clocked_on => CLK_port, Q => REGISTERS_3_8_port, QN => n_1119);
   REGISTERS_reg_3_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N175, next_state => N91, 
               clocked_on => CLK_port, Q => REGISTERS_3_7_port, QN => n_1120);
   REGISTERS_reg_3_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N175, next_state => N90, 
               clocked_on => CLK_port, Q => REGISTERS_3_6_port, QN => n_1121);
   REGISTERS_reg_3_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N175, next_state => N89, 
               clocked_on => CLK_port, Q => REGISTERS_3_5_port, QN => n_1122);
   REGISTERS_reg_3_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N175, next_state => N88, 
               clocked_on => CLK_port, Q => REGISTERS_3_4_port, QN => n_1123);
   REGISTERS_reg_3_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N175, next_state => N87, 
               clocked_on => CLK_port, Q => REGISTERS_3_3_port, QN => n_1124);
   REGISTERS_reg_3_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N175, next_state => N86, 
               clocked_on => CLK_port, Q => REGISTERS_3_2_port, QN => n_1125);
   REGISTERS_reg_3_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N175, next_state => N85, 
               clocked_on => CLK_port, Q => REGISTERS_3_1_port, QN => n_1126);
   REGISTERS_reg_3_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N175, next_state => N84, 
               clocked_on => CLK_port, Q => REGISTERS_3_0_port, QN => n_1127);
   REGISTERS_reg_4_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N174, next_state => N115, 
               clocked_on => CLK_port, Q => REGISTERS_4_31_port, QN => n_1128);
   REGISTERS_reg_4_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N174, next_state => N114, 
               clocked_on => CLK_port, Q => REGISTERS_4_30_port, QN => n_1129);
   REGISTERS_reg_4_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N174, next_state => N113, 
               clocked_on => CLK_port, Q => REGISTERS_4_29_port, QN => n_1130);
   REGISTERS_reg_4_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N174, next_state => N112, 
               clocked_on => CLK_port, Q => REGISTERS_4_28_port, QN => n_1131);
   REGISTERS_reg_4_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N174, next_state => N111, 
               clocked_on => CLK_port, Q => REGISTERS_4_27_port, QN => n_1132);
   REGISTERS_reg_4_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N174, next_state => N110, 
               clocked_on => CLK_port, Q => REGISTERS_4_26_port, QN => n_1133);
   REGISTERS_reg_4_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N174, next_state => N109, 
               clocked_on => CLK_port, Q => REGISTERS_4_25_port, QN => n_1134);
   REGISTERS_reg_4_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N174, next_state => N108, 
               clocked_on => CLK_port, Q => REGISTERS_4_24_port, QN => n_1135);
   REGISTERS_reg_4_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N174, next_state => N107, 
               clocked_on => CLK_port, Q => REGISTERS_4_23_port, QN => n_1136);
   REGISTERS_reg_4_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N174, next_state => N106, 
               clocked_on => CLK_port, Q => REGISTERS_4_22_port, QN => n_1137);
   REGISTERS_reg_4_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N174, next_state => N105, 
               clocked_on => CLK_port, Q => REGISTERS_4_21_port, QN => n_1138);
   REGISTERS_reg_4_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N174, next_state => N104, 
               clocked_on => CLK_port, Q => REGISTERS_4_20_port, QN => n_1139);
   REGISTERS_reg_4_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N174, next_state => N103, 
               clocked_on => CLK_port, Q => REGISTERS_4_19_port, QN => n_1140);
   REGISTERS_reg_4_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N174, next_state => N102, 
               clocked_on => CLK_port, Q => REGISTERS_4_18_port, QN => n_1141);
   REGISTERS_reg_4_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N174, next_state => N101, 
               clocked_on => CLK_port, Q => REGISTERS_4_17_port, QN => n_1142);
   REGISTERS_reg_4_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N174, next_state => N100, 
               clocked_on => CLK_port, Q => REGISTERS_4_16_port, QN => n_1143);
   REGISTERS_reg_4_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N174, next_state => N99, 
               clocked_on => CLK_port, Q => REGISTERS_4_15_port, QN => n_1144);
   REGISTERS_reg_4_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N174, next_state => N98, 
               clocked_on => CLK_port, Q => REGISTERS_4_14_port, QN => n_1145);
   REGISTERS_reg_4_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N174, next_state => N97, 
               clocked_on => CLK_port, Q => REGISTERS_4_13_port, QN => n_1146);
   REGISTERS_reg_4_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N174, next_state => N96, 
               clocked_on => CLK_port, Q => REGISTERS_4_12_port, QN => n_1147);
   REGISTERS_reg_4_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N174, next_state => N95, 
               clocked_on => CLK_port, Q => REGISTERS_4_11_port, QN => n_1148);
   REGISTERS_reg_4_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N174, next_state => N94, 
               clocked_on => CLK_port, Q => REGISTERS_4_10_port, QN => n_1149);
   REGISTERS_reg_4_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N174, next_state => N93, 
               clocked_on => CLK_port, Q => REGISTERS_4_9_port, QN => n_1150);
   REGISTERS_reg_4_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N174, next_state => N92, 
               clocked_on => CLK_port, Q => REGISTERS_4_8_port, QN => n_1151);
   REGISTERS_reg_4_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N174, next_state => N91, 
               clocked_on => CLK_port, Q => REGISTERS_4_7_port, QN => n_1152);
   REGISTERS_reg_4_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N174, next_state => N90, 
               clocked_on => CLK_port, Q => REGISTERS_4_6_port, QN => n_1153);
   REGISTERS_reg_4_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N174, next_state => N89, 
               clocked_on => CLK_port, Q => REGISTERS_4_5_port, QN => n_1154);
   REGISTERS_reg_4_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N174, next_state => N88, 
               clocked_on => CLK_port, Q => REGISTERS_4_4_port, QN => n_1155);
   REGISTERS_reg_4_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N174, next_state => N87, 
               clocked_on => CLK_port, Q => REGISTERS_4_3_port, QN => n_1156);
   REGISTERS_reg_4_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N174, next_state => N86, 
               clocked_on => CLK_port, Q => REGISTERS_4_2_port, QN => n_1157);
   REGISTERS_reg_4_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N174, next_state => N85, 
               clocked_on => CLK_port, Q => REGISTERS_4_1_port, QN => n_1158);
   REGISTERS_reg_4_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N174, next_state => N84, 
               clocked_on => CLK_port, Q => REGISTERS_4_0_port, QN => n_1159);
   REGISTERS_reg_5_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N173, next_state => N115, 
               clocked_on => CLK_port, Q => REGISTERS_5_31_port, QN => n_1160);
   REGISTERS_reg_5_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N173, next_state => N114, 
               clocked_on => CLK_port, Q => REGISTERS_5_30_port, QN => n_1161);
   REGISTERS_reg_5_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N173, next_state => N113, 
               clocked_on => CLK_port, Q => REGISTERS_5_29_port, QN => n_1162);
   REGISTERS_reg_5_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N173, next_state => N112, 
               clocked_on => CLK_port, Q => REGISTERS_5_28_port, QN => n_1163);
   REGISTERS_reg_5_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N173, next_state => N111, 
               clocked_on => CLK_port, Q => REGISTERS_5_27_port, QN => n_1164);
   REGISTERS_reg_5_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N173, next_state => N110, 
               clocked_on => CLK_port, Q => REGISTERS_5_26_port, QN => n_1165);
   REGISTERS_reg_5_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N173, next_state => N109, 
               clocked_on => CLK_port, Q => REGISTERS_5_25_port, QN => n_1166);
   REGISTERS_reg_5_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N173, next_state => N108, 
               clocked_on => CLK_port, Q => REGISTERS_5_24_port, QN => n_1167);
   REGISTERS_reg_5_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N173, next_state => N107, 
               clocked_on => CLK_port, Q => REGISTERS_5_23_port, QN => n_1168);
   REGISTERS_reg_5_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N173, next_state => N106, 
               clocked_on => CLK_port, Q => REGISTERS_5_22_port, QN => n_1169);
   REGISTERS_reg_5_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N173, next_state => N105, 
               clocked_on => CLK_port, Q => REGISTERS_5_21_port, QN => n_1170);
   REGISTERS_reg_5_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N173, next_state => N104, 
               clocked_on => CLK_port, Q => REGISTERS_5_20_port, QN => n_1171);
   REGISTERS_reg_5_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N173, next_state => N103, 
               clocked_on => CLK_port, Q => REGISTERS_5_19_port, QN => n_1172);
   REGISTERS_reg_5_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N173, next_state => N102, 
               clocked_on => CLK_port, Q => REGISTERS_5_18_port, QN => n_1173);
   REGISTERS_reg_5_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N173, next_state => N101, 
               clocked_on => CLK_port, Q => REGISTERS_5_17_port, QN => n_1174);
   REGISTERS_reg_5_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N173, next_state => N100, 
               clocked_on => CLK_port, Q => REGISTERS_5_16_port, QN => n_1175);
   REGISTERS_reg_5_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N173, next_state => N99, 
               clocked_on => CLK_port, Q => REGISTERS_5_15_port, QN => n_1176);
   REGISTERS_reg_5_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N173, next_state => N98, 
               clocked_on => CLK_port, Q => REGISTERS_5_14_port, QN => n_1177);
   REGISTERS_reg_5_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N173, next_state => N97, 
               clocked_on => CLK_port, Q => REGISTERS_5_13_port, QN => n_1178);
   REGISTERS_reg_5_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N173, next_state => N96, 
               clocked_on => CLK_port, Q => REGISTERS_5_12_port, QN => n_1179);
   REGISTERS_reg_5_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N173, next_state => N95, 
               clocked_on => CLK_port, Q => REGISTERS_5_11_port, QN => n_1180);
   REGISTERS_reg_5_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N173, next_state => N94, 
               clocked_on => CLK_port, Q => REGISTERS_5_10_port, QN => n_1181);
   REGISTERS_reg_5_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N173, next_state => N93, 
               clocked_on => CLK_port, Q => REGISTERS_5_9_port, QN => n_1182);
   REGISTERS_reg_5_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N173, next_state => N92, 
               clocked_on => CLK_port, Q => REGISTERS_5_8_port, QN => n_1183);
   REGISTERS_reg_5_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N173, next_state => N91, 
               clocked_on => CLK_port, Q => REGISTERS_5_7_port, QN => n_1184);
   REGISTERS_reg_5_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N173, next_state => N90, 
               clocked_on => CLK_port, Q => REGISTERS_5_6_port, QN => n_1185);
   REGISTERS_reg_5_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N173, next_state => N89, 
               clocked_on => CLK_port, Q => REGISTERS_5_5_port, QN => n_1186);
   REGISTERS_reg_5_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N173, next_state => N88, 
               clocked_on => CLK_port, Q => REGISTERS_5_4_port, QN => n_1187);
   REGISTERS_reg_5_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N173, next_state => N87, 
               clocked_on => CLK_port, Q => REGISTERS_5_3_port, QN => n_1188);
   REGISTERS_reg_5_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N173, next_state => N86, 
               clocked_on => CLK_port, Q => REGISTERS_5_2_port, QN => n_1189);
   REGISTERS_reg_5_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N173, next_state => N85, 
               clocked_on => CLK_port, Q => REGISTERS_5_1_port, QN => n_1190);
   REGISTERS_reg_5_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N173, next_state => N84, 
               clocked_on => CLK_port, Q => REGISTERS_5_0_port, QN => n_1191);
   REGISTERS_reg_6_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N172, next_state => N115, 
               clocked_on => CLK_port, Q => REGISTERS_6_31_port, QN => n_1192);
   REGISTERS_reg_6_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N172, next_state => N114, 
               clocked_on => CLK_port, Q => REGISTERS_6_30_port, QN => n_1193);
   REGISTERS_reg_6_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N172, next_state => N113, 
               clocked_on => CLK_port, Q => REGISTERS_6_29_port, QN => n_1194);
   REGISTERS_reg_6_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N172, next_state => N112, 
               clocked_on => CLK_port, Q => REGISTERS_6_28_port, QN => n_1195);
   REGISTERS_reg_6_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N172, next_state => N111, 
               clocked_on => CLK_port, Q => REGISTERS_6_27_port, QN => n_1196);
   REGISTERS_reg_6_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N172, next_state => N110, 
               clocked_on => CLK_port, Q => REGISTERS_6_26_port, QN => n_1197);
   REGISTERS_reg_6_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N172, next_state => N109, 
               clocked_on => CLK_port, Q => REGISTERS_6_25_port, QN => n_1198);
   REGISTERS_reg_6_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N172, next_state => N108, 
               clocked_on => CLK_port, Q => REGISTERS_6_24_port, QN => n_1199);
   REGISTERS_reg_6_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N172, next_state => N107, 
               clocked_on => CLK_port, Q => REGISTERS_6_23_port, QN => n_1200);
   REGISTERS_reg_6_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N172, next_state => N106, 
               clocked_on => CLK_port, Q => REGISTERS_6_22_port, QN => n_1201);
   REGISTERS_reg_6_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N172, next_state => N105, 
               clocked_on => CLK_port, Q => REGISTERS_6_21_port, QN => n_1202);
   REGISTERS_reg_6_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N172, next_state => N104, 
               clocked_on => CLK_port, Q => REGISTERS_6_20_port, QN => n_1203);
   REGISTERS_reg_6_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N172, next_state => N103, 
               clocked_on => CLK_port, Q => REGISTERS_6_19_port, QN => n_1204);
   REGISTERS_reg_6_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N172, next_state => N102, 
               clocked_on => CLK_port, Q => REGISTERS_6_18_port, QN => n_1205);
   REGISTERS_reg_6_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N172, next_state => N101, 
               clocked_on => CLK_port, Q => REGISTERS_6_17_port, QN => n_1206);
   REGISTERS_reg_6_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N172, next_state => N100, 
               clocked_on => CLK_port, Q => REGISTERS_6_16_port, QN => n_1207);
   REGISTERS_reg_6_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N172, next_state => N99, 
               clocked_on => CLK_port, Q => REGISTERS_6_15_port, QN => n_1208);
   REGISTERS_reg_6_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N172, next_state => N98, 
               clocked_on => CLK_port, Q => REGISTERS_6_14_port, QN => n_1209);
   REGISTERS_reg_6_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N172, next_state => N97, 
               clocked_on => CLK_port, Q => REGISTERS_6_13_port, QN => n_1210);
   REGISTERS_reg_6_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N172, next_state => N96, 
               clocked_on => CLK_port, Q => REGISTERS_6_12_port, QN => n_1211);
   REGISTERS_reg_6_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N172, next_state => N95, 
               clocked_on => CLK_port, Q => REGISTERS_6_11_port, QN => n_1212);
   REGISTERS_reg_6_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N172, next_state => N94, 
               clocked_on => CLK_port, Q => REGISTERS_6_10_port, QN => n_1213);
   REGISTERS_reg_6_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N172, next_state => N93, 
               clocked_on => CLK_port, Q => REGISTERS_6_9_port, QN => n_1214);
   REGISTERS_reg_6_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N172, next_state => N92, 
               clocked_on => CLK_port, Q => REGISTERS_6_8_port, QN => n_1215);
   REGISTERS_reg_6_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N172, next_state => N91, 
               clocked_on => CLK_port, Q => REGISTERS_6_7_port, QN => n_1216);
   REGISTERS_reg_6_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N172, next_state => N90, 
               clocked_on => CLK_port, Q => REGISTERS_6_6_port, QN => n_1217);
   REGISTERS_reg_6_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N172, next_state => N89, 
               clocked_on => CLK_port, Q => REGISTERS_6_5_port, QN => n_1218);
   REGISTERS_reg_6_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N172, next_state => N88, 
               clocked_on => CLK_port, Q => REGISTERS_6_4_port, QN => n_1219);
   REGISTERS_reg_6_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N172, next_state => N87, 
               clocked_on => CLK_port, Q => REGISTERS_6_3_port, QN => n_1220);
   REGISTERS_reg_6_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N172, next_state => N86, 
               clocked_on => CLK_port, Q => REGISTERS_6_2_port, QN => n_1221);
   REGISTERS_reg_6_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N172, next_state => N85, 
               clocked_on => CLK_port, Q => REGISTERS_6_1_port, QN => n_1222);
   REGISTERS_reg_6_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N172, next_state => N84, 
               clocked_on => CLK_port, Q => REGISTERS_6_0_port, QN => n_1223);
   REGISTERS_reg_7_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N171, next_state => N115, 
               clocked_on => CLK_port, Q => REGISTERS_7_31_port, QN => n_1224);
   REGISTERS_reg_7_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N171, next_state => N114, 
               clocked_on => CLK_port, Q => REGISTERS_7_30_port, QN => n_1225);
   REGISTERS_reg_7_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N171, next_state => N113, 
               clocked_on => CLK_port, Q => REGISTERS_7_29_port, QN => n_1226);
   REGISTERS_reg_7_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N171, next_state => N112, 
               clocked_on => CLK_port, Q => REGISTERS_7_28_port, QN => n_1227);
   REGISTERS_reg_7_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N171, next_state => N111, 
               clocked_on => CLK_port, Q => REGISTERS_7_27_port, QN => n_1228);
   REGISTERS_reg_7_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N171, next_state => N110, 
               clocked_on => CLK_port, Q => REGISTERS_7_26_port, QN => n_1229);
   REGISTERS_reg_7_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N171, next_state => N109, 
               clocked_on => CLK_port, Q => REGISTERS_7_25_port, QN => n_1230);
   REGISTERS_reg_7_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N171, next_state => N108, 
               clocked_on => CLK_port, Q => REGISTERS_7_24_port, QN => n_1231);
   REGISTERS_reg_7_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N171, next_state => N107, 
               clocked_on => CLK_port, Q => REGISTERS_7_23_port, QN => n_1232);
   REGISTERS_reg_7_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N171, next_state => N106, 
               clocked_on => CLK_port, Q => REGISTERS_7_22_port, QN => n_1233);
   REGISTERS_reg_7_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N171, next_state => N105, 
               clocked_on => CLK_port, Q => REGISTERS_7_21_port, QN => n_1234);
   REGISTERS_reg_7_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N171, next_state => N104, 
               clocked_on => CLK_port, Q => REGISTERS_7_20_port, QN => n_1235);
   REGISTERS_reg_7_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N171, next_state => N103, 
               clocked_on => CLK_port, Q => REGISTERS_7_19_port, QN => n_1236);
   REGISTERS_reg_7_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N171, next_state => N102, 
               clocked_on => CLK_port, Q => REGISTERS_7_18_port, QN => n_1237);
   REGISTERS_reg_7_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N171, next_state => N101, 
               clocked_on => CLK_port, Q => REGISTERS_7_17_port, QN => n_1238);
   REGISTERS_reg_7_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N171, next_state => N100, 
               clocked_on => CLK_port, Q => REGISTERS_7_16_port, QN => n_1239);
   REGISTERS_reg_7_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N171, next_state => N99, 
               clocked_on => CLK_port, Q => REGISTERS_7_15_port, QN => n_1240);
   REGISTERS_reg_7_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N171, next_state => N98, 
               clocked_on => CLK_port, Q => REGISTERS_7_14_port, QN => n_1241);
   REGISTERS_reg_7_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N171, next_state => N97, 
               clocked_on => CLK_port, Q => REGISTERS_7_13_port, QN => n_1242);
   REGISTERS_reg_7_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N171, next_state => N96, 
               clocked_on => CLK_port, Q => REGISTERS_7_12_port, QN => n_1243);
   REGISTERS_reg_7_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N171, next_state => N95, 
               clocked_on => CLK_port, Q => REGISTERS_7_11_port, QN => n_1244);
   REGISTERS_reg_7_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N171, next_state => N94, 
               clocked_on => CLK_port, Q => REGISTERS_7_10_port, QN => n_1245);
   REGISTERS_reg_7_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N171, next_state => N93, 
               clocked_on => CLK_port, Q => REGISTERS_7_9_port, QN => n_1246);
   REGISTERS_reg_7_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N171, next_state => N92, 
               clocked_on => CLK_port, Q => REGISTERS_7_8_port, QN => n_1247);
   REGISTERS_reg_7_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N171, next_state => N91, 
               clocked_on => CLK_port, Q => REGISTERS_7_7_port, QN => n_1248);
   REGISTERS_reg_7_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N171, next_state => N90, 
               clocked_on => CLK_port, Q => REGISTERS_7_6_port, QN => n_1249);
   REGISTERS_reg_7_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N171, next_state => N89, 
               clocked_on => CLK_port, Q => REGISTERS_7_5_port, QN => n_1250);
   REGISTERS_reg_7_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N171, next_state => N88, 
               clocked_on => CLK_port, Q => REGISTERS_7_4_port, QN => n_1251);
   REGISTERS_reg_7_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N171, next_state => N87, 
               clocked_on => CLK_port, Q => REGISTERS_7_3_port, QN => n_1252);
   REGISTERS_reg_7_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N171, next_state => N86, 
               clocked_on => CLK_port, Q => REGISTERS_7_2_port, QN => n_1253);
   REGISTERS_reg_7_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N171, next_state => N85, 
               clocked_on => CLK_port, Q => REGISTERS_7_1_port, QN => n_1254);
   REGISTERS_reg_7_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N171, next_state => N84, 
               clocked_on => CLK_port, Q => REGISTERS_7_0_port, QN => n_1255);
   REGISTERS_reg_8_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N170, next_state => N115, 
               clocked_on => CLK_port, Q => REGISTERS_8_31_port, QN => n_1256);
   REGISTERS_reg_8_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N170, next_state => N114, 
               clocked_on => CLK_port, Q => REGISTERS_8_30_port, QN => n_1257);
   REGISTERS_reg_8_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N170, next_state => N113, 
               clocked_on => CLK_port, Q => REGISTERS_8_29_port, QN => n_1258);
   REGISTERS_reg_8_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N170, next_state => N112, 
               clocked_on => CLK_port, Q => REGISTERS_8_28_port, QN => n_1259);
   REGISTERS_reg_8_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N170, next_state => N111, 
               clocked_on => CLK_port, Q => REGISTERS_8_27_port, QN => n_1260);
   REGISTERS_reg_8_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N170, next_state => N110, 
               clocked_on => CLK_port, Q => REGISTERS_8_26_port, QN => n_1261);
   REGISTERS_reg_8_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N170, next_state => N109, 
               clocked_on => CLK_port, Q => REGISTERS_8_25_port, QN => n_1262);
   REGISTERS_reg_8_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N170, next_state => N108, 
               clocked_on => CLK_port, Q => REGISTERS_8_24_port, QN => n_1263);
   REGISTERS_reg_8_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N170, next_state => N107, 
               clocked_on => CLK_port, Q => REGISTERS_8_23_port, QN => n_1264);
   REGISTERS_reg_8_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N170, next_state => N106, 
               clocked_on => CLK_port, Q => REGISTERS_8_22_port, QN => n_1265);
   REGISTERS_reg_8_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N170, next_state => N105, 
               clocked_on => CLK_port, Q => REGISTERS_8_21_port, QN => n_1266);
   REGISTERS_reg_8_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N170, next_state => N104, 
               clocked_on => CLK_port, Q => REGISTERS_8_20_port, QN => n_1267);
   REGISTERS_reg_8_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N170, next_state => N103, 
               clocked_on => CLK_port, Q => REGISTERS_8_19_port, QN => n_1268);
   REGISTERS_reg_8_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N170, next_state => N102, 
               clocked_on => CLK_port, Q => REGISTERS_8_18_port, QN => n_1269);
   REGISTERS_reg_8_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N170, next_state => N101, 
               clocked_on => CLK_port, Q => REGISTERS_8_17_port, QN => n_1270);
   REGISTERS_reg_8_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N170, next_state => N100, 
               clocked_on => CLK_port, Q => REGISTERS_8_16_port, QN => n_1271);
   REGISTERS_reg_8_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N170, next_state => N99, 
               clocked_on => CLK_port, Q => REGISTERS_8_15_port, QN => n_1272);
   REGISTERS_reg_8_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N170, next_state => N98, 
               clocked_on => CLK_port, Q => REGISTERS_8_14_port, QN => n_1273);
   REGISTERS_reg_8_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N170, next_state => N97, 
               clocked_on => CLK_port, Q => REGISTERS_8_13_port, QN => n_1274);
   REGISTERS_reg_8_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N170, next_state => N96, 
               clocked_on => CLK_port, Q => REGISTERS_8_12_port, QN => n_1275);
   REGISTERS_reg_8_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N170, next_state => N95, 
               clocked_on => CLK_port, Q => REGISTERS_8_11_port, QN => n_1276);
   REGISTERS_reg_8_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N170, next_state => N94, 
               clocked_on => CLK_port, Q => REGISTERS_8_10_port, QN => n_1277);
   REGISTERS_reg_8_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N170, next_state => N93, 
               clocked_on => CLK_port, Q => REGISTERS_8_9_port, QN => n_1278);
   REGISTERS_reg_8_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N170, next_state => N92, 
               clocked_on => CLK_port, Q => REGISTERS_8_8_port, QN => n_1279);
   REGISTERS_reg_8_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N170, next_state => N91, 
               clocked_on => CLK_port, Q => REGISTERS_8_7_port, QN => n_1280);
   REGISTERS_reg_8_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N170, next_state => N90, 
               clocked_on => CLK_port, Q => REGISTERS_8_6_port, QN => n_1281);
   REGISTERS_reg_8_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N170, next_state => N89, 
               clocked_on => CLK_port, Q => REGISTERS_8_5_port, QN => n_1282);
   REGISTERS_reg_8_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N170, next_state => N88, 
               clocked_on => CLK_port, Q => REGISTERS_8_4_port, QN => n_1283);
   REGISTERS_reg_8_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N170, next_state => N87, 
               clocked_on => CLK_port, Q => REGISTERS_8_3_port, QN => n_1284);
   REGISTERS_reg_8_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N170, next_state => N86, 
               clocked_on => CLK_port, Q => REGISTERS_8_2_port, QN => n_1285);
   REGISTERS_reg_8_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N170, next_state => N85, 
               clocked_on => CLK_port, Q => REGISTERS_8_1_port, QN => n_1286);
   REGISTERS_reg_8_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N170, next_state => N84, 
               clocked_on => CLK_port, Q => REGISTERS_8_0_port, QN => n_1287);
   REGISTERS_reg_9_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N169, next_state => N115, 
               clocked_on => CLK_port, Q => REGISTERS_9_31_port, QN => n_1288);
   REGISTERS_reg_9_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N169, next_state => N114, 
               clocked_on => CLK_port, Q => REGISTERS_9_30_port, QN => n_1289);
   REGISTERS_reg_9_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N169, next_state => N113, 
               clocked_on => CLK_port, Q => REGISTERS_9_29_port, QN => n_1290);
   REGISTERS_reg_9_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N169, next_state => N112, 
               clocked_on => CLK_port, Q => REGISTERS_9_28_port, QN => n_1291);
   REGISTERS_reg_9_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N169, next_state => N111, 
               clocked_on => CLK_port, Q => REGISTERS_9_27_port, QN => n_1292);
   REGISTERS_reg_9_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N169, next_state => N110, 
               clocked_on => CLK_port, Q => REGISTERS_9_26_port, QN => n_1293);
   REGISTERS_reg_9_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N169, next_state => N109, 
               clocked_on => CLK_port, Q => REGISTERS_9_25_port, QN => n_1294);
   REGISTERS_reg_9_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N169, next_state => N108, 
               clocked_on => CLK_port, Q => REGISTERS_9_24_port, QN => n_1295);
   REGISTERS_reg_9_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N169, next_state => N107, 
               clocked_on => CLK_port, Q => REGISTERS_9_23_port, QN => n_1296);
   REGISTERS_reg_9_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N169, next_state => N106, 
               clocked_on => CLK_port, Q => REGISTERS_9_22_port, QN => n_1297);
   REGISTERS_reg_9_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N169, next_state => N105, 
               clocked_on => CLK_port, Q => REGISTERS_9_21_port, QN => n_1298);
   REGISTERS_reg_9_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N169, next_state => N104, 
               clocked_on => CLK_port, Q => REGISTERS_9_20_port, QN => n_1299);
   REGISTERS_reg_9_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N169, next_state => N103, 
               clocked_on => CLK_port, Q => REGISTERS_9_19_port, QN => n_1300);
   REGISTERS_reg_9_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N169, next_state => N102, 
               clocked_on => CLK_port, Q => REGISTERS_9_18_port, QN => n_1301);
   REGISTERS_reg_9_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N169, next_state => N101, 
               clocked_on => CLK_port, Q => REGISTERS_9_17_port, QN => n_1302);
   REGISTERS_reg_9_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N169, next_state => N100, 
               clocked_on => CLK_port, Q => REGISTERS_9_16_port, QN => n_1303);
   REGISTERS_reg_9_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N169, next_state => N99, 
               clocked_on => CLK_port, Q => REGISTERS_9_15_port, QN => n_1304);
   REGISTERS_reg_9_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N169, next_state => N98, 
               clocked_on => CLK_port, Q => REGISTERS_9_14_port, QN => n_1305);
   REGISTERS_reg_9_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N169, next_state => N97, 
               clocked_on => CLK_port, Q => REGISTERS_9_13_port, QN => n_1306);
   REGISTERS_reg_9_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N169, next_state => N96, 
               clocked_on => CLK_port, Q => REGISTERS_9_12_port, QN => n_1307);
   REGISTERS_reg_9_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N169, next_state => N95, 
               clocked_on => CLK_port, Q => REGISTERS_9_11_port, QN => n_1308);
   REGISTERS_reg_9_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N169, next_state => N94, 
               clocked_on => CLK_port, Q => REGISTERS_9_10_port, QN => n_1309);
   REGISTERS_reg_9_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N169, next_state => N93, 
               clocked_on => CLK_port, Q => REGISTERS_9_9_port, QN => n_1310);
   REGISTERS_reg_9_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N169, next_state => N92, 
               clocked_on => CLK_port, Q => REGISTERS_9_8_port, QN => n_1311);
   REGISTERS_reg_9_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N169, next_state => N91, 
               clocked_on => CLK_port, Q => REGISTERS_9_7_port, QN => n_1312);
   REGISTERS_reg_9_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N169, next_state => N90, 
               clocked_on => CLK_port, Q => REGISTERS_9_6_port, QN => n_1313);
   REGISTERS_reg_9_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N169, next_state => N89, 
               clocked_on => CLK_port, Q => REGISTERS_9_5_port, QN => n_1314);
   REGISTERS_reg_9_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N169, next_state => N88, 
               clocked_on => CLK_port, Q => REGISTERS_9_4_port, QN => n_1315);
   REGISTERS_reg_9_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N169, next_state => N87, 
               clocked_on => CLK_port, Q => REGISTERS_9_3_port, QN => n_1316);
   REGISTERS_reg_9_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N169, next_state => N86, 
               clocked_on => CLK_port, Q => REGISTERS_9_2_port, QN => n_1317);
   REGISTERS_reg_9_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N169, next_state => N85, 
               clocked_on => CLK_port, Q => REGISTERS_9_1_port, QN => n_1318);
   REGISTERS_reg_9_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N169, next_state => N84, 
               clocked_on => CLK_port, Q => REGISTERS_9_0_port, QN => n_1319);
   REGISTERS_reg_10_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N168, next_state => N115, 
               clocked_on => CLK_port, Q => REGISTERS_10_31_port, QN => n_1320
               );
   REGISTERS_reg_10_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N168, next_state => N114, 
               clocked_on => CLK_port, Q => REGISTERS_10_30_port, QN => n_1321
               );
   REGISTERS_reg_10_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N168, next_state => N113, 
               clocked_on => CLK_port, Q => REGISTERS_10_29_port, QN => n_1322
               );
   REGISTERS_reg_10_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N168, next_state => N112, 
               clocked_on => CLK_port, Q => REGISTERS_10_28_port, QN => n_1323
               );
   REGISTERS_reg_10_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N168, next_state => N111, 
               clocked_on => CLK_port, Q => REGISTERS_10_27_port, QN => n_1324
               );
   REGISTERS_reg_10_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N168, next_state => N110, 
               clocked_on => CLK_port, Q => REGISTERS_10_26_port, QN => n_1325
               );
   REGISTERS_reg_10_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N168, next_state => N109, 
               clocked_on => CLK_port, Q => REGISTERS_10_25_port, QN => n_1326
               );
   REGISTERS_reg_10_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N168, next_state => N108, 
               clocked_on => CLK_port, Q => REGISTERS_10_24_port, QN => n_1327
               );
   REGISTERS_reg_10_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N168, next_state => N107, 
               clocked_on => CLK_port, Q => REGISTERS_10_23_port, QN => n_1328
               );
   REGISTERS_reg_10_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N168, next_state => N106, 
               clocked_on => CLK_port, Q => REGISTERS_10_22_port, QN => n_1329
               );
   REGISTERS_reg_10_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N168, next_state => N105, 
               clocked_on => CLK_port, Q => REGISTERS_10_21_port, QN => n_1330
               );
   REGISTERS_reg_10_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N168, next_state => N104, 
               clocked_on => CLK_port, Q => REGISTERS_10_20_port, QN => n_1331
               );
   REGISTERS_reg_10_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N168, next_state => N103, 
               clocked_on => CLK_port, Q => REGISTERS_10_19_port, QN => n_1332
               );
   REGISTERS_reg_10_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N168, next_state => N102, 
               clocked_on => CLK_port, Q => REGISTERS_10_18_port, QN => n_1333
               );
   REGISTERS_reg_10_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N168, next_state => N101, 
               clocked_on => CLK_port, Q => REGISTERS_10_17_port, QN => n_1334
               );
   REGISTERS_reg_10_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N168, next_state => N100, 
               clocked_on => CLK_port, Q => REGISTERS_10_16_port, QN => n_1335
               );
   REGISTERS_reg_10_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N168, next_state => N99, 
               clocked_on => CLK_port, Q => REGISTERS_10_15_port, QN => n_1336
               );
   REGISTERS_reg_10_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N168, next_state => N98, 
               clocked_on => CLK_port, Q => REGISTERS_10_14_port, QN => n_1337
               );
   REGISTERS_reg_10_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N168, next_state => N97, 
               clocked_on => CLK_port, Q => REGISTERS_10_13_port, QN => n_1338
               );
   REGISTERS_reg_10_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N168, next_state => N96, 
               clocked_on => CLK_port, Q => REGISTERS_10_12_port, QN => n_1339
               );
   REGISTERS_reg_10_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N168, next_state => N95, 
               clocked_on => CLK_port, Q => REGISTERS_10_11_port, QN => n_1340
               );
   REGISTERS_reg_10_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N168, next_state => N94, 
               clocked_on => CLK_port, Q => REGISTERS_10_10_port, QN => n_1341
               );
   REGISTERS_reg_10_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N168, next_state => N93, 
               clocked_on => CLK_port, Q => REGISTERS_10_9_port, QN => n_1342);
   REGISTERS_reg_10_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N168, next_state => N92, 
               clocked_on => CLK_port, Q => REGISTERS_10_8_port, QN => n_1343);
   REGISTERS_reg_10_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N168, next_state => N91, 
               clocked_on => CLK_port, Q => REGISTERS_10_7_port, QN => n_1344);
   REGISTERS_reg_10_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N168, next_state => N90, 
               clocked_on => CLK_port, Q => REGISTERS_10_6_port, QN => n_1345);
   REGISTERS_reg_10_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N168, next_state => N89, 
               clocked_on => CLK_port, Q => REGISTERS_10_5_port, QN => n_1346);
   REGISTERS_reg_10_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N168, next_state => N88, 
               clocked_on => CLK_port, Q => REGISTERS_10_4_port, QN => n_1347);
   REGISTERS_reg_10_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N168, next_state => N87, 
               clocked_on => CLK_port, Q => REGISTERS_10_3_port, QN => n_1348);
   REGISTERS_reg_10_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N168, next_state => N86, 
               clocked_on => CLK_port, Q => REGISTERS_10_2_port, QN => n_1349);
   REGISTERS_reg_10_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N168, next_state => N85, 
               clocked_on => CLK_port, Q => REGISTERS_10_1_port, QN => n_1350);
   REGISTERS_reg_10_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N168, next_state => N84, 
               clocked_on => CLK_port, Q => REGISTERS_10_0_port, QN => n_1351);
   REGISTERS_reg_11_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N167, next_state => N115, 
               clocked_on => CLK_port, Q => REGISTERS_11_31_port, QN => n_1352
               );
   REGISTERS_reg_11_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N167, next_state => N114, 
               clocked_on => CLK_port, Q => REGISTERS_11_30_port, QN => n_1353
               );
   REGISTERS_reg_11_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N167, next_state => N113, 
               clocked_on => CLK_port, Q => REGISTERS_11_29_port, QN => n_1354
               );
   REGISTERS_reg_11_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N167, next_state => N112, 
               clocked_on => CLK_port, Q => REGISTERS_11_28_port, QN => n_1355
               );
   REGISTERS_reg_11_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N167, next_state => N111, 
               clocked_on => CLK_port, Q => REGISTERS_11_27_port, QN => n_1356
               );
   REGISTERS_reg_11_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N167, next_state => N110, 
               clocked_on => CLK_port, Q => REGISTERS_11_26_port, QN => n_1357
               );
   REGISTERS_reg_11_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N167, next_state => N109, 
               clocked_on => CLK_port, Q => REGISTERS_11_25_port, QN => n_1358
               );
   REGISTERS_reg_11_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N167, next_state => N108, 
               clocked_on => CLK_port, Q => REGISTERS_11_24_port, QN => n_1359
               );
   REGISTERS_reg_11_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N167, next_state => N107, 
               clocked_on => CLK_port, Q => REGISTERS_11_23_port, QN => n_1360
               );
   REGISTERS_reg_11_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N167, next_state => N106, 
               clocked_on => CLK_port, Q => REGISTERS_11_22_port, QN => n_1361
               );
   REGISTERS_reg_11_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N167, next_state => N105, 
               clocked_on => CLK_port, Q => REGISTERS_11_21_port, QN => n_1362
               );
   REGISTERS_reg_11_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N167, next_state => N104, 
               clocked_on => CLK_port, Q => REGISTERS_11_20_port, QN => n_1363
               );
   REGISTERS_reg_11_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N167, next_state => N103, 
               clocked_on => CLK_port, Q => REGISTERS_11_19_port, QN => n_1364
               );
   REGISTERS_reg_11_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N167, next_state => N102, 
               clocked_on => CLK_port, Q => REGISTERS_11_18_port, QN => n_1365
               );
   REGISTERS_reg_11_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N167, next_state => N101, 
               clocked_on => CLK_port, Q => REGISTERS_11_17_port, QN => n_1366
               );
   REGISTERS_reg_11_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N167, next_state => N100, 
               clocked_on => CLK_port, Q => REGISTERS_11_16_port, QN => n_1367
               );
   REGISTERS_reg_11_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N167, next_state => N99, 
               clocked_on => CLK_port, Q => REGISTERS_11_15_port, QN => n_1368
               );
   REGISTERS_reg_11_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N167, next_state => N98, 
               clocked_on => CLK_port, Q => REGISTERS_11_14_port, QN => n_1369
               );
   REGISTERS_reg_11_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N167, next_state => N97, 
               clocked_on => CLK_port, Q => REGISTERS_11_13_port, QN => n_1370
               );
   REGISTERS_reg_11_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N167, next_state => N96, 
               clocked_on => CLK_port, Q => REGISTERS_11_12_port, QN => n_1371
               );
   REGISTERS_reg_11_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N167, next_state => N95, 
               clocked_on => CLK_port, Q => REGISTERS_11_11_port, QN => n_1372
               );
   REGISTERS_reg_11_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N167, next_state => N94, 
               clocked_on => CLK_port, Q => REGISTERS_11_10_port, QN => n_1373
               );
   REGISTERS_reg_11_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N167, next_state => N93, 
               clocked_on => CLK_port, Q => REGISTERS_11_9_port, QN => n_1374);
   REGISTERS_reg_11_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N167, next_state => N92, 
               clocked_on => CLK_port, Q => REGISTERS_11_8_port, QN => n_1375);
   REGISTERS_reg_11_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N167, next_state => N91, 
               clocked_on => CLK_port, Q => REGISTERS_11_7_port, QN => n_1376);
   REGISTERS_reg_11_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N167, next_state => N90, 
               clocked_on => CLK_port, Q => REGISTERS_11_6_port, QN => n_1377);
   REGISTERS_reg_11_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N167, next_state => N89, 
               clocked_on => CLK_port, Q => REGISTERS_11_5_port, QN => n_1378);
   REGISTERS_reg_11_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N167, next_state => N88, 
               clocked_on => CLK_port, Q => REGISTERS_11_4_port, QN => n_1379);
   REGISTERS_reg_11_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N167, next_state => N87, 
               clocked_on => CLK_port, Q => REGISTERS_11_3_port, QN => n_1380);
   REGISTERS_reg_11_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N167, next_state => N86, 
               clocked_on => CLK_port, Q => REGISTERS_11_2_port, QN => n_1381);
   REGISTERS_reg_11_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N167, next_state => N85, 
               clocked_on => CLK_port, Q => REGISTERS_11_1_port, QN => n_1382);
   REGISTERS_reg_11_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N167, next_state => N84, 
               clocked_on => CLK_port, Q => REGISTERS_11_0_port, QN => n_1383);
   REGISTERS_reg_12_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N166, next_state => N115, 
               clocked_on => CLK_port, Q => REGISTERS_12_31_port, QN => n_1384
               );
   REGISTERS_reg_12_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N166, next_state => N114, 
               clocked_on => CLK_port, Q => REGISTERS_12_30_port, QN => n_1385
               );
   REGISTERS_reg_12_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N166, next_state => N113, 
               clocked_on => CLK_port, Q => REGISTERS_12_29_port, QN => n_1386
               );
   REGISTERS_reg_12_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N166, next_state => N112, 
               clocked_on => CLK_port, Q => REGISTERS_12_28_port, QN => n_1387
               );
   REGISTERS_reg_12_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N166, next_state => N111, 
               clocked_on => CLK_port, Q => REGISTERS_12_27_port, QN => n_1388
               );
   REGISTERS_reg_12_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N166, next_state => N110, 
               clocked_on => CLK_port, Q => REGISTERS_12_26_port, QN => n_1389
               );
   REGISTERS_reg_12_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N166, next_state => N109, 
               clocked_on => CLK_port, Q => REGISTERS_12_25_port, QN => n_1390
               );
   REGISTERS_reg_12_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N166, next_state => N108, 
               clocked_on => CLK_port, Q => REGISTERS_12_24_port, QN => n_1391
               );
   REGISTERS_reg_12_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N166, next_state => N107, 
               clocked_on => CLK_port, Q => REGISTERS_12_23_port, QN => n_1392
               );
   REGISTERS_reg_12_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N166, next_state => N106, 
               clocked_on => CLK_port, Q => REGISTERS_12_22_port, QN => n_1393
               );
   REGISTERS_reg_12_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N166, next_state => N105, 
               clocked_on => CLK_port, Q => REGISTERS_12_21_port, QN => n_1394
               );
   REGISTERS_reg_12_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N166, next_state => N104, 
               clocked_on => CLK_port, Q => REGISTERS_12_20_port, QN => n_1395
               );
   REGISTERS_reg_12_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N166, next_state => N103, 
               clocked_on => CLK_port, Q => REGISTERS_12_19_port, QN => n_1396
               );
   REGISTERS_reg_12_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N166, next_state => N102, 
               clocked_on => CLK_port, Q => REGISTERS_12_18_port, QN => n_1397
               );
   REGISTERS_reg_12_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N166, next_state => N101, 
               clocked_on => CLK_port, Q => REGISTERS_12_17_port, QN => n_1398
               );
   REGISTERS_reg_12_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N166, next_state => N100, 
               clocked_on => CLK_port, Q => REGISTERS_12_16_port, QN => n_1399
               );
   REGISTERS_reg_12_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N166, next_state => N99, 
               clocked_on => CLK_port, Q => REGISTERS_12_15_port, QN => n_1400
               );
   REGISTERS_reg_12_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N166, next_state => N98, 
               clocked_on => CLK_port, Q => REGISTERS_12_14_port, QN => n_1401
               );
   REGISTERS_reg_12_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N166, next_state => N97, 
               clocked_on => CLK_port, Q => REGISTERS_12_13_port, QN => n_1402
               );
   REGISTERS_reg_12_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N166, next_state => N96, 
               clocked_on => CLK_port, Q => REGISTERS_12_12_port, QN => n_1403
               );
   REGISTERS_reg_12_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N166, next_state => N95, 
               clocked_on => CLK_port, Q => REGISTERS_12_11_port, QN => n_1404
               );
   REGISTERS_reg_12_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N166, next_state => N94, 
               clocked_on => CLK_port, Q => REGISTERS_12_10_port, QN => n_1405
               );
   REGISTERS_reg_12_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N166, next_state => N93, 
               clocked_on => CLK_port, Q => REGISTERS_12_9_port, QN => n_1406);
   REGISTERS_reg_12_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N166, next_state => N92, 
               clocked_on => CLK_port, Q => REGISTERS_12_8_port, QN => n_1407);
   REGISTERS_reg_12_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N166, next_state => N91, 
               clocked_on => CLK_port, Q => REGISTERS_12_7_port, QN => n_1408);
   REGISTERS_reg_12_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N166, next_state => N90, 
               clocked_on => CLK_port, Q => REGISTERS_12_6_port, QN => n_1409);
   REGISTERS_reg_12_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N166, next_state => N89, 
               clocked_on => CLK_port, Q => REGISTERS_12_5_port, QN => n_1410);
   REGISTERS_reg_12_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N166, next_state => N88, 
               clocked_on => CLK_port, Q => REGISTERS_12_4_port, QN => n_1411);
   REGISTERS_reg_12_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N166, next_state => N87, 
               clocked_on => CLK_port, Q => REGISTERS_12_3_port, QN => n_1412);
   REGISTERS_reg_12_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N166, next_state => N86, 
               clocked_on => CLK_port, Q => REGISTERS_12_2_port, QN => n_1413);
   REGISTERS_reg_12_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N166, next_state => N85, 
               clocked_on => CLK_port, Q => REGISTERS_12_1_port, QN => n_1414);
   REGISTERS_reg_12_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N166, next_state => N84, 
               clocked_on => CLK_port, Q => REGISTERS_12_0_port, QN => n_1415);
   REGISTERS_reg_13_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N165, next_state => N115, 
               clocked_on => CLK_port, Q => REGISTERS_13_31_port, QN => n_1416
               );
   REGISTERS_reg_13_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N165, next_state => N114, 
               clocked_on => CLK_port, Q => REGISTERS_13_30_port, QN => n_1417
               );
   REGISTERS_reg_13_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N165, next_state => N113, 
               clocked_on => CLK_port, Q => REGISTERS_13_29_port, QN => n_1418
               );
   REGISTERS_reg_13_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N165, next_state => N112, 
               clocked_on => CLK_port, Q => REGISTERS_13_28_port, QN => n_1419
               );
   REGISTERS_reg_13_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N165, next_state => N111, 
               clocked_on => CLK_port, Q => REGISTERS_13_27_port, QN => n_1420
               );
   REGISTERS_reg_13_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N165, next_state => N110, 
               clocked_on => CLK_port, Q => REGISTERS_13_26_port, QN => n_1421
               );
   REGISTERS_reg_13_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N165, next_state => N109, 
               clocked_on => CLK_port, Q => REGISTERS_13_25_port, QN => n_1422
               );
   REGISTERS_reg_13_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N165, next_state => N108, 
               clocked_on => CLK_port, Q => REGISTERS_13_24_port, QN => n_1423
               );
   REGISTERS_reg_13_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N165, next_state => N107, 
               clocked_on => CLK_port, Q => REGISTERS_13_23_port, QN => n_1424
               );
   REGISTERS_reg_13_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N165, next_state => N106, 
               clocked_on => CLK_port, Q => REGISTERS_13_22_port, QN => n_1425
               );
   REGISTERS_reg_13_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N165, next_state => N105, 
               clocked_on => CLK_port, Q => REGISTERS_13_21_port, QN => n_1426
               );
   REGISTERS_reg_13_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N165, next_state => N104, 
               clocked_on => CLK_port, Q => REGISTERS_13_20_port, QN => n_1427
               );
   REGISTERS_reg_13_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N165, next_state => N103, 
               clocked_on => CLK_port, Q => REGISTERS_13_19_port, QN => n_1428
               );
   REGISTERS_reg_13_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N165, next_state => N102, 
               clocked_on => CLK_port, Q => REGISTERS_13_18_port, QN => n_1429
               );
   REGISTERS_reg_13_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N165, next_state => N101, 
               clocked_on => CLK_port, Q => REGISTERS_13_17_port, QN => n_1430
               );
   REGISTERS_reg_13_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N165, next_state => N100, 
               clocked_on => CLK_port, Q => REGISTERS_13_16_port, QN => n_1431
               );
   REGISTERS_reg_13_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N165, next_state => N99, 
               clocked_on => CLK_port, Q => REGISTERS_13_15_port, QN => n_1432
               );
   REGISTERS_reg_13_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N165, next_state => N98, 
               clocked_on => CLK_port, Q => REGISTERS_13_14_port, QN => n_1433
               );
   REGISTERS_reg_13_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N165, next_state => N97, 
               clocked_on => CLK_port, Q => REGISTERS_13_13_port, QN => n_1434
               );
   REGISTERS_reg_13_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N165, next_state => N96, 
               clocked_on => CLK_port, Q => REGISTERS_13_12_port, QN => n_1435
               );
   REGISTERS_reg_13_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N165, next_state => N95, 
               clocked_on => CLK_port, Q => REGISTERS_13_11_port, QN => n_1436
               );
   REGISTERS_reg_13_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N165, next_state => N94, 
               clocked_on => CLK_port, Q => REGISTERS_13_10_port, QN => n_1437
               );
   REGISTERS_reg_13_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N165, next_state => N93, 
               clocked_on => CLK_port, Q => REGISTERS_13_9_port, QN => n_1438);
   REGISTERS_reg_13_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N165, next_state => N92, 
               clocked_on => CLK_port, Q => REGISTERS_13_8_port, QN => n_1439);
   REGISTERS_reg_13_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N165, next_state => N91, 
               clocked_on => CLK_port, Q => REGISTERS_13_7_port, QN => n_1440);
   REGISTERS_reg_13_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N165, next_state => N90, 
               clocked_on => CLK_port, Q => REGISTERS_13_6_port, QN => n_1441);
   REGISTERS_reg_13_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N165, next_state => N89, 
               clocked_on => CLK_port, Q => REGISTERS_13_5_port, QN => n_1442);
   REGISTERS_reg_13_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N165, next_state => N88, 
               clocked_on => CLK_port, Q => REGISTERS_13_4_port, QN => n_1443);
   REGISTERS_reg_13_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N165, next_state => N87, 
               clocked_on => CLK_port, Q => REGISTERS_13_3_port, QN => n_1444);
   REGISTERS_reg_13_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N165, next_state => N86, 
               clocked_on => CLK_port, Q => REGISTERS_13_2_port, QN => n_1445);
   REGISTERS_reg_13_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N165, next_state => N85, 
               clocked_on => CLK_port, Q => REGISTERS_13_1_port, QN => n_1446);
   REGISTERS_reg_13_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N165, next_state => N84, 
               clocked_on => CLK_port, Q => REGISTERS_13_0_port, QN => n_1447);
   REGISTERS_reg_14_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N164, next_state => N115, 
               clocked_on => CLK_port, Q => REGISTERS_14_31_port, QN => n_1448
               );
   REGISTERS_reg_14_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N164, next_state => N114, 
               clocked_on => CLK_port, Q => REGISTERS_14_30_port, QN => n_1449
               );
   REGISTERS_reg_14_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N164, next_state => N113, 
               clocked_on => CLK_port, Q => REGISTERS_14_29_port, QN => n_1450
               );
   REGISTERS_reg_14_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N164, next_state => N112, 
               clocked_on => CLK_port, Q => REGISTERS_14_28_port, QN => n_1451
               );
   REGISTERS_reg_14_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N164, next_state => N111, 
               clocked_on => CLK_port, Q => REGISTERS_14_27_port, QN => n_1452
               );
   REGISTERS_reg_14_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N164, next_state => N110, 
               clocked_on => CLK_port, Q => REGISTERS_14_26_port, QN => n_1453
               );
   REGISTERS_reg_14_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N164, next_state => N109, 
               clocked_on => CLK_port, Q => REGISTERS_14_25_port, QN => n_1454
               );
   REGISTERS_reg_14_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N164, next_state => N108, 
               clocked_on => CLK_port, Q => REGISTERS_14_24_port, QN => n_1455
               );
   REGISTERS_reg_14_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N164, next_state => N107, 
               clocked_on => CLK_port, Q => REGISTERS_14_23_port, QN => n_1456
               );
   REGISTERS_reg_14_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N164, next_state => N106, 
               clocked_on => CLK_port, Q => REGISTERS_14_22_port, QN => n_1457
               );
   REGISTERS_reg_14_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N164, next_state => N105, 
               clocked_on => CLK_port, Q => REGISTERS_14_21_port, QN => n_1458
               );
   REGISTERS_reg_14_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N164, next_state => N104, 
               clocked_on => CLK_port, Q => REGISTERS_14_20_port, QN => n_1459
               );
   REGISTERS_reg_14_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N164, next_state => N103, 
               clocked_on => CLK_port, Q => REGISTERS_14_19_port, QN => n_1460
               );
   REGISTERS_reg_14_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N164, next_state => N102, 
               clocked_on => CLK_port, Q => REGISTERS_14_18_port, QN => n_1461
               );
   REGISTERS_reg_14_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N164, next_state => N101, 
               clocked_on => CLK_port, Q => REGISTERS_14_17_port, QN => n_1462
               );
   REGISTERS_reg_14_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N164, next_state => N100, 
               clocked_on => CLK_port, Q => REGISTERS_14_16_port, QN => n_1463
               );
   REGISTERS_reg_14_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N164, next_state => N99, 
               clocked_on => CLK_port, Q => REGISTERS_14_15_port, QN => n_1464
               );
   REGISTERS_reg_14_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N164, next_state => N98, 
               clocked_on => CLK_port, Q => REGISTERS_14_14_port, QN => n_1465
               );
   REGISTERS_reg_14_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N164, next_state => N97, 
               clocked_on => CLK_port, Q => REGISTERS_14_13_port, QN => n_1466
               );
   REGISTERS_reg_14_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N164, next_state => N96, 
               clocked_on => CLK_port, Q => REGISTERS_14_12_port, QN => n_1467
               );
   REGISTERS_reg_14_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N164, next_state => N95, 
               clocked_on => CLK_port, Q => REGISTERS_14_11_port, QN => n_1468
               );
   REGISTERS_reg_14_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N164, next_state => N94, 
               clocked_on => CLK_port, Q => REGISTERS_14_10_port, QN => n_1469
               );
   REGISTERS_reg_14_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N164, next_state => N93, 
               clocked_on => CLK_port, Q => REGISTERS_14_9_port, QN => n_1470);
   REGISTERS_reg_14_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N164, next_state => N92, 
               clocked_on => CLK_port, Q => REGISTERS_14_8_port, QN => n_1471);
   REGISTERS_reg_14_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N164, next_state => N91, 
               clocked_on => CLK_port, Q => REGISTERS_14_7_port, QN => n_1472);
   REGISTERS_reg_14_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N164, next_state => N90, 
               clocked_on => CLK_port, Q => REGISTERS_14_6_port, QN => n_1473);
   REGISTERS_reg_14_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N164, next_state => N89, 
               clocked_on => CLK_port, Q => REGISTERS_14_5_port, QN => n_1474);
   REGISTERS_reg_14_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N164, next_state => N88, 
               clocked_on => CLK_port, Q => REGISTERS_14_4_port, QN => n_1475);
   REGISTERS_reg_14_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N164, next_state => N87, 
               clocked_on => CLK_port, Q => REGISTERS_14_3_port, QN => n_1476);
   REGISTERS_reg_14_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N164, next_state => N86, 
               clocked_on => CLK_port, Q => REGISTERS_14_2_port, QN => n_1477);
   REGISTERS_reg_14_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N164, next_state => N85, 
               clocked_on => CLK_port, Q => REGISTERS_14_1_port, QN => n_1478);
   REGISTERS_reg_14_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N164, next_state => N84, 
               clocked_on => CLK_port, Q => REGISTERS_14_0_port, QN => n_1479);
   REGISTERS_reg_15_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N163, next_state => N115, 
               clocked_on => CLK_port, Q => REGISTERS_15_31_port, QN => n_1480
               );
   REGISTERS_reg_15_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N163, next_state => N114, 
               clocked_on => CLK_port, Q => REGISTERS_15_30_port, QN => n_1481
               );
   REGISTERS_reg_15_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N163, next_state => N113, 
               clocked_on => CLK_port, Q => REGISTERS_15_29_port, QN => n_1482
               );
   REGISTERS_reg_15_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N163, next_state => N112, 
               clocked_on => CLK_port, Q => REGISTERS_15_28_port, QN => n_1483
               );
   REGISTERS_reg_15_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N163, next_state => N111, 
               clocked_on => CLK_port, Q => REGISTERS_15_27_port, QN => n_1484
               );
   REGISTERS_reg_15_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N163, next_state => N110, 
               clocked_on => CLK_port, Q => REGISTERS_15_26_port, QN => n_1485
               );
   REGISTERS_reg_15_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N163, next_state => N109, 
               clocked_on => CLK_port, Q => REGISTERS_15_25_port, QN => n_1486
               );
   REGISTERS_reg_15_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N163, next_state => N108, 
               clocked_on => CLK_port, Q => REGISTERS_15_24_port, QN => n_1487
               );
   REGISTERS_reg_15_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N163, next_state => N107, 
               clocked_on => CLK_port, Q => REGISTERS_15_23_port, QN => n_1488
               );
   REGISTERS_reg_15_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N163, next_state => N106, 
               clocked_on => CLK_port, Q => REGISTERS_15_22_port, QN => n_1489
               );
   REGISTERS_reg_15_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N163, next_state => N105, 
               clocked_on => CLK_port, Q => REGISTERS_15_21_port, QN => n_1490
               );
   REGISTERS_reg_15_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N163, next_state => N104, 
               clocked_on => CLK_port, Q => REGISTERS_15_20_port, QN => n_1491
               );
   REGISTERS_reg_15_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N163, next_state => N103, 
               clocked_on => CLK_port, Q => REGISTERS_15_19_port, QN => n_1492
               );
   REGISTERS_reg_15_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N163, next_state => N102, 
               clocked_on => CLK_port, Q => REGISTERS_15_18_port, QN => n_1493
               );
   REGISTERS_reg_15_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N163, next_state => N101, 
               clocked_on => CLK_port, Q => REGISTERS_15_17_port, QN => n_1494
               );
   REGISTERS_reg_15_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N163, next_state => N100, 
               clocked_on => CLK_port, Q => REGISTERS_15_16_port, QN => n_1495
               );
   REGISTERS_reg_15_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N163, next_state => N99, 
               clocked_on => CLK_port, Q => REGISTERS_15_15_port, QN => n_1496
               );
   REGISTERS_reg_15_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N163, next_state => N98, 
               clocked_on => CLK_port, Q => REGISTERS_15_14_port, QN => n_1497
               );
   REGISTERS_reg_15_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N163, next_state => N97, 
               clocked_on => CLK_port, Q => REGISTERS_15_13_port, QN => n_1498
               );
   REGISTERS_reg_15_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N163, next_state => N96, 
               clocked_on => CLK_port, Q => REGISTERS_15_12_port, QN => n_1499
               );
   REGISTERS_reg_15_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N163, next_state => N95, 
               clocked_on => CLK_port, Q => REGISTERS_15_11_port, QN => n_1500
               );
   REGISTERS_reg_15_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N163, next_state => N94, 
               clocked_on => CLK_port, Q => REGISTERS_15_10_port, QN => n_1501
               );
   REGISTERS_reg_15_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N163, next_state => N93, 
               clocked_on => CLK_port, Q => REGISTERS_15_9_port, QN => n_1502);
   REGISTERS_reg_15_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N163, next_state => N92, 
               clocked_on => CLK_port, Q => REGISTERS_15_8_port, QN => n_1503);
   REGISTERS_reg_15_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N163, next_state => N91, 
               clocked_on => CLK_port, Q => REGISTERS_15_7_port, QN => n_1504);
   REGISTERS_reg_15_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N163, next_state => N90, 
               clocked_on => CLK_port, Q => REGISTERS_15_6_port, QN => n_1505);
   REGISTERS_reg_15_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N163, next_state => N89, 
               clocked_on => CLK_port, Q => REGISTERS_15_5_port, QN => n_1506);
   REGISTERS_reg_15_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N163, next_state => N88, 
               clocked_on => CLK_port, Q => REGISTERS_15_4_port, QN => n_1507);
   REGISTERS_reg_15_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N163, next_state => N87, 
               clocked_on => CLK_port, Q => REGISTERS_15_3_port, QN => n_1508);
   REGISTERS_reg_15_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N163, next_state => N86, 
               clocked_on => CLK_port, Q => REGISTERS_15_2_port, QN => n_1509);
   REGISTERS_reg_15_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N163, next_state => N85, 
               clocked_on => CLK_port, Q => REGISTERS_15_1_port, QN => n_1510);
   REGISTERS_reg_15_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N163, next_state => N84, 
               clocked_on => CLK_port, Q => REGISTERS_15_0_port, QN => n_1511);
   REGISTERS_reg_16_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N162, next_state => N115, 
               clocked_on => CLK_port, Q => REGISTERS_16_31_port, QN => n_1512
               );
   REGISTERS_reg_16_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N162, next_state => N114, 
               clocked_on => CLK_port, Q => REGISTERS_16_30_port, QN => n_1513
               );
   REGISTERS_reg_16_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N162, next_state => N113, 
               clocked_on => CLK_port, Q => REGISTERS_16_29_port, QN => n_1514
               );
   REGISTERS_reg_16_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N162, next_state => N112, 
               clocked_on => CLK_port, Q => REGISTERS_16_28_port, QN => n_1515
               );
   REGISTERS_reg_16_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N162, next_state => N111, 
               clocked_on => CLK_port, Q => REGISTERS_16_27_port, QN => n_1516
               );
   REGISTERS_reg_16_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N162, next_state => N110, 
               clocked_on => CLK_port, Q => REGISTERS_16_26_port, QN => n_1517
               );
   REGISTERS_reg_16_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N162, next_state => N109, 
               clocked_on => CLK_port, Q => REGISTERS_16_25_port, QN => n_1518
               );
   REGISTERS_reg_16_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N162, next_state => N108, 
               clocked_on => CLK_port, Q => REGISTERS_16_24_port, QN => n_1519
               );
   REGISTERS_reg_16_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N162, next_state => N107, 
               clocked_on => CLK_port, Q => REGISTERS_16_23_port, QN => n_1520
               );
   REGISTERS_reg_16_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N162, next_state => N106, 
               clocked_on => CLK_port, Q => REGISTERS_16_22_port, QN => n_1521
               );
   REGISTERS_reg_16_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N162, next_state => N105, 
               clocked_on => CLK_port, Q => REGISTERS_16_21_port, QN => n_1522
               );
   REGISTERS_reg_16_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N162, next_state => N104, 
               clocked_on => CLK_port, Q => REGISTERS_16_20_port, QN => n_1523
               );
   REGISTERS_reg_16_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N162, next_state => N103, 
               clocked_on => CLK_port, Q => REGISTERS_16_19_port, QN => n_1524
               );
   REGISTERS_reg_16_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N162, next_state => N102, 
               clocked_on => CLK_port, Q => REGISTERS_16_18_port, QN => n_1525
               );
   REGISTERS_reg_16_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N162, next_state => N101, 
               clocked_on => CLK_port, Q => REGISTERS_16_17_port, QN => n_1526
               );
   REGISTERS_reg_16_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N162, next_state => N100, 
               clocked_on => CLK_port, Q => REGISTERS_16_16_port, QN => n_1527
               );
   REGISTERS_reg_16_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N162, next_state => N99, 
               clocked_on => CLK_port, Q => REGISTERS_16_15_port, QN => n_1528
               );
   REGISTERS_reg_16_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N162, next_state => N98, 
               clocked_on => CLK_port, Q => REGISTERS_16_14_port, QN => n_1529
               );
   REGISTERS_reg_16_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N162, next_state => N97, 
               clocked_on => CLK_port, Q => REGISTERS_16_13_port, QN => n_1530
               );
   REGISTERS_reg_16_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N162, next_state => N96, 
               clocked_on => CLK_port, Q => REGISTERS_16_12_port, QN => n_1531
               );
   REGISTERS_reg_16_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N162, next_state => N95, 
               clocked_on => CLK_port, Q => REGISTERS_16_11_port, QN => n_1532
               );
   REGISTERS_reg_16_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N162, next_state => N94, 
               clocked_on => CLK_port, Q => REGISTERS_16_10_port, QN => n_1533
               );
   REGISTERS_reg_16_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N162, next_state => N93, 
               clocked_on => CLK_port, Q => REGISTERS_16_9_port, QN => n_1534);
   REGISTERS_reg_16_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N162, next_state => N92, 
               clocked_on => CLK_port, Q => REGISTERS_16_8_port, QN => n_1535);
   REGISTERS_reg_16_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N162, next_state => N91, 
               clocked_on => CLK_port, Q => REGISTERS_16_7_port, QN => n_1536);
   REGISTERS_reg_16_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N162, next_state => N90, 
               clocked_on => CLK_port, Q => REGISTERS_16_6_port, QN => n_1537);
   REGISTERS_reg_16_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N162, next_state => N89, 
               clocked_on => CLK_port, Q => REGISTERS_16_5_port, QN => n_1538);
   REGISTERS_reg_16_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N162, next_state => N88, 
               clocked_on => CLK_port, Q => REGISTERS_16_4_port, QN => n_1539);
   REGISTERS_reg_16_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N162, next_state => N87, 
               clocked_on => CLK_port, Q => REGISTERS_16_3_port, QN => n_1540);
   REGISTERS_reg_16_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N162, next_state => N86, 
               clocked_on => CLK_port, Q => REGISTERS_16_2_port, QN => n_1541);
   REGISTERS_reg_16_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N162, next_state => N85, 
               clocked_on => CLK_port, Q => REGISTERS_16_1_port, QN => n_1542);
   REGISTERS_reg_16_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N162, next_state => N84, 
               clocked_on => CLK_port, Q => REGISTERS_16_0_port, QN => n_1543);
   REGISTERS_reg_17_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N161, next_state => N115, 
               clocked_on => CLK_port, Q => REGISTERS_17_31_port, QN => n_1544
               );
   REGISTERS_reg_17_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N161, next_state => N114, 
               clocked_on => CLK_port, Q => REGISTERS_17_30_port, QN => n_1545
               );
   REGISTERS_reg_17_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N161, next_state => N113, 
               clocked_on => CLK_port, Q => REGISTERS_17_29_port, QN => n_1546
               );
   REGISTERS_reg_17_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N161, next_state => N112, 
               clocked_on => CLK_port, Q => REGISTERS_17_28_port, QN => n_1547
               );
   REGISTERS_reg_17_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N161, next_state => N111, 
               clocked_on => CLK_port, Q => REGISTERS_17_27_port, QN => n_1548
               );
   REGISTERS_reg_17_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N161, next_state => N110, 
               clocked_on => CLK_port, Q => REGISTERS_17_26_port, QN => n_1549
               );
   REGISTERS_reg_17_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N161, next_state => N109, 
               clocked_on => CLK_port, Q => REGISTERS_17_25_port, QN => n_1550
               );
   REGISTERS_reg_17_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N161, next_state => N108, 
               clocked_on => CLK_port, Q => REGISTERS_17_24_port, QN => n_1551
               );
   REGISTERS_reg_17_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N161, next_state => N107, 
               clocked_on => CLK_port, Q => REGISTERS_17_23_port, QN => n_1552
               );
   REGISTERS_reg_17_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N161, next_state => N106, 
               clocked_on => CLK_port, Q => REGISTERS_17_22_port, QN => n_1553
               );
   REGISTERS_reg_17_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N161, next_state => N105, 
               clocked_on => CLK_port, Q => REGISTERS_17_21_port, QN => n_1554
               );
   REGISTERS_reg_17_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N161, next_state => N104, 
               clocked_on => CLK_port, Q => REGISTERS_17_20_port, QN => n_1555
               );
   REGISTERS_reg_17_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N161, next_state => N103, 
               clocked_on => CLK_port, Q => REGISTERS_17_19_port, QN => n_1556
               );
   REGISTERS_reg_17_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N161, next_state => N102, 
               clocked_on => CLK_port, Q => REGISTERS_17_18_port, QN => n_1557
               );
   REGISTERS_reg_17_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N161, next_state => N101, 
               clocked_on => CLK_port, Q => REGISTERS_17_17_port, QN => n_1558
               );
   REGISTERS_reg_17_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N161, next_state => N100, 
               clocked_on => CLK_port, Q => REGISTERS_17_16_port, QN => n_1559
               );
   REGISTERS_reg_17_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N161, next_state => N99, 
               clocked_on => CLK_port, Q => REGISTERS_17_15_port, QN => n_1560
               );
   REGISTERS_reg_17_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N161, next_state => N98, 
               clocked_on => CLK_port, Q => REGISTERS_17_14_port, QN => n_1561
               );
   REGISTERS_reg_17_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N161, next_state => N97, 
               clocked_on => CLK_port, Q => REGISTERS_17_13_port, QN => n_1562
               );
   REGISTERS_reg_17_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N161, next_state => N96, 
               clocked_on => CLK_port, Q => REGISTERS_17_12_port, QN => n_1563
               );
   REGISTERS_reg_17_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N161, next_state => N95, 
               clocked_on => CLK_port, Q => REGISTERS_17_11_port, QN => n_1564
               );
   REGISTERS_reg_17_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N161, next_state => N94, 
               clocked_on => CLK_port, Q => REGISTERS_17_10_port, QN => n_1565
               );
   REGISTERS_reg_17_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N161, next_state => N93, 
               clocked_on => CLK_port, Q => REGISTERS_17_9_port, QN => n_1566);
   REGISTERS_reg_17_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N161, next_state => N92, 
               clocked_on => CLK_port, Q => REGISTERS_17_8_port, QN => n_1567);
   REGISTERS_reg_17_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N161, next_state => N91, 
               clocked_on => CLK_port, Q => REGISTERS_17_7_port, QN => n_1568);
   REGISTERS_reg_17_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N161, next_state => N90, 
               clocked_on => CLK_port, Q => REGISTERS_17_6_port, QN => n_1569);
   REGISTERS_reg_17_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N161, next_state => N89, 
               clocked_on => CLK_port, Q => REGISTERS_17_5_port, QN => n_1570);
   REGISTERS_reg_17_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N161, next_state => N88, 
               clocked_on => CLK_port, Q => REGISTERS_17_4_port, QN => n_1571);
   REGISTERS_reg_17_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N161, next_state => N87, 
               clocked_on => CLK_port, Q => REGISTERS_17_3_port, QN => n_1572);
   REGISTERS_reg_17_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N161, next_state => N86, 
               clocked_on => CLK_port, Q => REGISTERS_17_2_port, QN => n_1573);
   REGISTERS_reg_17_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N161, next_state => N85, 
               clocked_on => CLK_port, Q => REGISTERS_17_1_port, QN => n_1574);
   REGISTERS_reg_17_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N161, next_state => N84, 
               clocked_on => CLK_port, Q => REGISTERS_17_0_port, QN => n_1575);
   REGISTERS_reg_18_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N160, next_state => N115, 
               clocked_on => CLK_port, Q => REGISTERS_18_31_port, QN => n_1576
               );
   REGISTERS_reg_18_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N160, next_state => N114, 
               clocked_on => CLK_port, Q => REGISTERS_18_30_port, QN => n_1577
               );
   REGISTERS_reg_18_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N160, next_state => N113, 
               clocked_on => CLK_port, Q => REGISTERS_18_29_port, QN => n_1578
               );
   REGISTERS_reg_18_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N160, next_state => N112, 
               clocked_on => CLK_port, Q => REGISTERS_18_28_port, QN => n_1579
               );
   REGISTERS_reg_18_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N160, next_state => N111, 
               clocked_on => CLK_port, Q => REGISTERS_18_27_port, QN => n_1580
               );
   REGISTERS_reg_18_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N160, next_state => N110, 
               clocked_on => CLK_port, Q => REGISTERS_18_26_port, QN => n_1581
               );
   REGISTERS_reg_18_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N160, next_state => N109, 
               clocked_on => CLK_port, Q => REGISTERS_18_25_port, QN => n_1582
               );
   REGISTERS_reg_18_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N160, next_state => N108, 
               clocked_on => CLK_port, Q => REGISTERS_18_24_port, QN => n_1583
               );
   REGISTERS_reg_18_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N160, next_state => N107, 
               clocked_on => CLK_port, Q => REGISTERS_18_23_port, QN => n_1584
               );
   REGISTERS_reg_18_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N160, next_state => N106, 
               clocked_on => CLK_port, Q => REGISTERS_18_22_port, QN => n_1585
               );
   REGISTERS_reg_18_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N160, next_state => N105, 
               clocked_on => CLK_port, Q => REGISTERS_18_21_port, QN => n_1586
               );
   REGISTERS_reg_18_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N160, next_state => N104, 
               clocked_on => CLK_port, Q => REGISTERS_18_20_port, QN => n_1587
               );
   REGISTERS_reg_18_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N160, next_state => N103, 
               clocked_on => CLK_port, Q => REGISTERS_18_19_port, QN => n_1588
               );
   REGISTERS_reg_18_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N160, next_state => N102, 
               clocked_on => CLK_port, Q => REGISTERS_18_18_port, QN => n_1589
               );
   REGISTERS_reg_18_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N160, next_state => N101, 
               clocked_on => CLK_port, Q => REGISTERS_18_17_port, QN => n_1590
               );
   REGISTERS_reg_18_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N160, next_state => N100, 
               clocked_on => CLK_port, Q => REGISTERS_18_16_port, QN => n_1591
               );
   REGISTERS_reg_18_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N160, next_state => N99, 
               clocked_on => CLK_port, Q => REGISTERS_18_15_port, QN => n_1592
               );
   REGISTERS_reg_18_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N160, next_state => N98, 
               clocked_on => CLK_port, Q => REGISTERS_18_14_port, QN => n_1593
               );
   REGISTERS_reg_18_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N160, next_state => N97, 
               clocked_on => CLK_port, Q => REGISTERS_18_13_port, QN => n_1594
               );
   REGISTERS_reg_18_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N160, next_state => N96, 
               clocked_on => CLK_port, Q => REGISTERS_18_12_port, QN => n_1595
               );
   REGISTERS_reg_18_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N160, next_state => N95, 
               clocked_on => CLK_port, Q => REGISTERS_18_11_port, QN => n_1596
               );
   REGISTERS_reg_18_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N160, next_state => N94, 
               clocked_on => CLK_port, Q => REGISTERS_18_10_port, QN => n_1597
               );
   REGISTERS_reg_18_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N160, next_state => N93, 
               clocked_on => CLK_port, Q => REGISTERS_18_9_port, QN => n_1598);
   REGISTERS_reg_18_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N160, next_state => N92, 
               clocked_on => CLK_port, Q => REGISTERS_18_8_port, QN => n_1599);
   REGISTERS_reg_18_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N160, next_state => N91, 
               clocked_on => CLK_port, Q => REGISTERS_18_7_port, QN => n_1600);
   REGISTERS_reg_18_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N160, next_state => N90, 
               clocked_on => CLK_port, Q => REGISTERS_18_6_port, QN => n_1601);
   REGISTERS_reg_18_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N160, next_state => N89, 
               clocked_on => CLK_port, Q => REGISTERS_18_5_port, QN => n_1602);
   REGISTERS_reg_18_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N160, next_state => N88, 
               clocked_on => CLK_port, Q => REGISTERS_18_4_port, QN => n_1603);
   REGISTERS_reg_18_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N160, next_state => N87, 
               clocked_on => CLK_port, Q => REGISTERS_18_3_port, QN => n_1604);
   REGISTERS_reg_18_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N160, next_state => N86, 
               clocked_on => CLK_port, Q => REGISTERS_18_2_port, QN => n_1605);
   REGISTERS_reg_18_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N160, next_state => N85, 
               clocked_on => CLK_port, Q => REGISTERS_18_1_port, QN => n_1606);
   REGISTERS_reg_18_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N160, next_state => N84, 
               clocked_on => CLK_port, Q => REGISTERS_18_0_port, QN => n_1607);
   REGISTERS_reg_19_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N159, next_state => N115, 
               clocked_on => CLK_port, Q => REGISTERS_19_31_port, QN => n_1608
               );
   REGISTERS_reg_19_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N159, next_state => N114, 
               clocked_on => CLK_port, Q => REGISTERS_19_30_port, QN => n_1609
               );
   REGISTERS_reg_19_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N159, next_state => N113, 
               clocked_on => CLK_port, Q => REGISTERS_19_29_port, QN => n_1610
               );
   REGISTERS_reg_19_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N159, next_state => N112, 
               clocked_on => CLK_port, Q => REGISTERS_19_28_port, QN => n_1611
               );
   REGISTERS_reg_19_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N159, next_state => N111, 
               clocked_on => CLK_port, Q => REGISTERS_19_27_port, QN => n_1612
               );
   REGISTERS_reg_19_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N159, next_state => N110, 
               clocked_on => CLK_port, Q => REGISTERS_19_26_port, QN => n_1613
               );
   REGISTERS_reg_19_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N159, next_state => N109, 
               clocked_on => CLK_port, Q => REGISTERS_19_25_port, QN => n_1614
               );
   REGISTERS_reg_19_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N159, next_state => N108, 
               clocked_on => CLK_port, Q => REGISTERS_19_24_port, QN => n_1615
               );
   REGISTERS_reg_19_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N159, next_state => N107, 
               clocked_on => CLK_port, Q => REGISTERS_19_23_port, QN => n_1616
               );
   REGISTERS_reg_19_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N159, next_state => N106, 
               clocked_on => CLK_port, Q => REGISTERS_19_22_port, QN => n_1617
               );
   REGISTERS_reg_19_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N159, next_state => N105, 
               clocked_on => CLK_port, Q => REGISTERS_19_21_port, QN => n_1618
               );
   REGISTERS_reg_19_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N159, next_state => N104, 
               clocked_on => CLK_port, Q => REGISTERS_19_20_port, QN => n_1619
               );
   REGISTERS_reg_19_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N159, next_state => N103, 
               clocked_on => CLK_port, Q => REGISTERS_19_19_port, QN => n_1620
               );
   REGISTERS_reg_19_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N159, next_state => N102, 
               clocked_on => CLK_port, Q => REGISTERS_19_18_port, QN => n_1621
               );
   REGISTERS_reg_19_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N159, next_state => N101, 
               clocked_on => CLK_port, Q => REGISTERS_19_17_port, QN => n_1622
               );
   REGISTERS_reg_19_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N159, next_state => N100, 
               clocked_on => CLK_port, Q => REGISTERS_19_16_port, QN => n_1623
               );
   REGISTERS_reg_19_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N159, next_state => N99, 
               clocked_on => CLK_port, Q => REGISTERS_19_15_port, QN => n_1624
               );
   REGISTERS_reg_19_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N159, next_state => N98, 
               clocked_on => CLK_port, Q => REGISTERS_19_14_port, QN => n_1625
               );
   REGISTERS_reg_19_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N159, next_state => N97, 
               clocked_on => CLK_port, Q => REGISTERS_19_13_port, QN => n_1626
               );
   REGISTERS_reg_19_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N159, next_state => N96, 
               clocked_on => CLK_port, Q => REGISTERS_19_12_port, QN => n_1627
               );
   REGISTERS_reg_19_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N159, next_state => N95, 
               clocked_on => CLK_port, Q => REGISTERS_19_11_port, QN => n_1628
               );
   REGISTERS_reg_19_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N159, next_state => N94, 
               clocked_on => CLK_port, Q => REGISTERS_19_10_port, QN => n_1629
               );
   REGISTERS_reg_19_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N159, next_state => N93, 
               clocked_on => CLK_port, Q => REGISTERS_19_9_port, QN => n_1630);
   REGISTERS_reg_19_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N159, next_state => N92, 
               clocked_on => CLK_port, Q => REGISTERS_19_8_port, QN => n_1631);
   REGISTERS_reg_19_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N159, next_state => N91, 
               clocked_on => CLK_port, Q => REGISTERS_19_7_port, QN => n_1632);
   REGISTERS_reg_19_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N159, next_state => N90, 
               clocked_on => CLK_port, Q => REGISTERS_19_6_port, QN => n_1633);
   REGISTERS_reg_19_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N159, next_state => N89, 
               clocked_on => CLK_port, Q => REGISTERS_19_5_port, QN => n_1634);
   REGISTERS_reg_19_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N159, next_state => N88, 
               clocked_on => CLK_port, Q => REGISTERS_19_4_port, QN => n_1635);
   REGISTERS_reg_19_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N159, next_state => N87, 
               clocked_on => CLK_port, Q => REGISTERS_19_3_port, QN => n_1636);
   REGISTERS_reg_19_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N159, next_state => N86, 
               clocked_on => CLK_port, Q => REGISTERS_19_2_port, QN => n_1637);
   REGISTERS_reg_19_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N159, next_state => N85, 
               clocked_on => CLK_port, Q => REGISTERS_19_1_port, QN => n_1638);
   REGISTERS_reg_19_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N159, next_state => N84, 
               clocked_on => CLK_port, Q => REGISTERS_19_0_port, QN => n_1639);
   REGISTERS_reg_20_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N158, next_state => N115, 
               clocked_on => CLK_port, Q => REGISTERS_20_31_port, QN => n_1640
               );
   REGISTERS_reg_20_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N158, next_state => N114, 
               clocked_on => CLK_port, Q => REGISTERS_20_30_port, QN => n_1641
               );
   REGISTERS_reg_20_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N158, next_state => N113, 
               clocked_on => CLK_port, Q => REGISTERS_20_29_port, QN => n_1642
               );
   REGISTERS_reg_20_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N158, next_state => N112, 
               clocked_on => CLK_port, Q => REGISTERS_20_28_port, QN => n_1643
               );
   REGISTERS_reg_20_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N158, next_state => N111, 
               clocked_on => CLK_port, Q => REGISTERS_20_27_port, QN => n_1644
               );
   REGISTERS_reg_20_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N158, next_state => N110, 
               clocked_on => CLK_port, Q => REGISTERS_20_26_port, QN => n_1645
               );
   REGISTERS_reg_20_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N158, next_state => N109, 
               clocked_on => CLK_port, Q => REGISTERS_20_25_port, QN => n_1646
               );
   REGISTERS_reg_20_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N158, next_state => N108, 
               clocked_on => CLK_port, Q => REGISTERS_20_24_port, QN => n_1647
               );
   REGISTERS_reg_20_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N158, next_state => N107, 
               clocked_on => CLK_port, Q => REGISTERS_20_23_port, QN => n_1648
               );
   REGISTERS_reg_20_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N158, next_state => N106, 
               clocked_on => CLK_port, Q => REGISTERS_20_22_port, QN => n_1649
               );
   REGISTERS_reg_20_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N158, next_state => N105, 
               clocked_on => CLK_port, Q => REGISTERS_20_21_port, QN => n_1650
               );
   REGISTERS_reg_20_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N158, next_state => N104, 
               clocked_on => CLK_port, Q => REGISTERS_20_20_port, QN => n_1651
               );
   REGISTERS_reg_20_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N158, next_state => N103, 
               clocked_on => CLK_port, Q => REGISTERS_20_19_port, QN => n_1652
               );
   REGISTERS_reg_20_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N158, next_state => N102, 
               clocked_on => CLK_port, Q => REGISTERS_20_18_port, QN => n_1653
               );
   REGISTERS_reg_20_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N158, next_state => N101, 
               clocked_on => CLK_port, Q => REGISTERS_20_17_port, QN => n_1654
               );
   REGISTERS_reg_20_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N158, next_state => N100, 
               clocked_on => CLK_port, Q => REGISTERS_20_16_port, QN => n_1655
               );
   REGISTERS_reg_20_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N158, next_state => N99, 
               clocked_on => CLK_port, Q => REGISTERS_20_15_port, QN => n_1656
               );
   REGISTERS_reg_20_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N158, next_state => N98, 
               clocked_on => CLK_port, Q => REGISTERS_20_14_port, QN => n_1657
               );
   REGISTERS_reg_20_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N158, next_state => N97, 
               clocked_on => CLK_port, Q => REGISTERS_20_13_port, QN => n_1658
               );
   REGISTERS_reg_20_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N158, next_state => N96, 
               clocked_on => CLK_port, Q => REGISTERS_20_12_port, QN => n_1659
               );
   REGISTERS_reg_20_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N158, next_state => N95, 
               clocked_on => CLK_port, Q => REGISTERS_20_11_port, QN => n_1660
               );
   REGISTERS_reg_20_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N158, next_state => N94, 
               clocked_on => CLK_port, Q => REGISTERS_20_10_port, QN => n_1661
               );
   REGISTERS_reg_20_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N158, next_state => N93, 
               clocked_on => CLK_port, Q => REGISTERS_20_9_port, QN => n_1662);
   REGISTERS_reg_20_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N158, next_state => N92, 
               clocked_on => CLK_port, Q => REGISTERS_20_8_port, QN => n_1663);
   REGISTERS_reg_20_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N158, next_state => N91, 
               clocked_on => CLK_port, Q => REGISTERS_20_7_port, QN => n_1664);
   REGISTERS_reg_20_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N158, next_state => N90, 
               clocked_on => CLK_port, Q => REGISTERS_20_6_port, QN => n_1665);
   REGISTERS_reg_20_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N158, next_state => N89, 
               clocked_on => CLK_port, Q => REGISTERS_20_5_port, QN => n_1666);
   REGISTERS_reg_20_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N158, next_state => N88, 
               clocked_on => CLK_port, Q => REGISTERS_20_4_port, QN => n_1667);
   REGISTERS_reg_20_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N158, next_state => N87, 
               clocked_on => CLK_port, Q => REGISTERS_20_3_port, QN => n_1668);
   REGISTERS_reg_20_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N158, next_state => N86, 
               clocked_on => CLK_port, Q => REGISTERS_20_2_port, QN => n_1669);
   REGISTERS_reg_20_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N158, next_state => N85, 
               clocked_on => CLK_port, Q => REGISTERS_20_1_port, QN => n_1670);
   REGISTERS_reg_20_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N158, next_state => N84, 
               clocked_on => CLK_port, Q => REGISTERS_20_0_port, QN => n_1671);
   REGISTERS_reg_21_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N157, next_state => N115, 
               clocked_on => CLK_port, Q => REGISTERS_21_31_port, QN => n_1672
               );
   REGISTERS_reg_21_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N157, next_state => N114, 
               clocked_on => CLK_port, Q => REGISTERS_21_30_port, QN => n_1673
               );
   REGISTERS_reg_21_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N157, next_state => N113, 
               clocked_on => CLK_port, Q => REGISTERS_21_29_port, QN => n_1674
               );
   REGISTERS_reg_21_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N157, next_state => N112, 
               clocked_on => CLK_port, Q => REGISTERS_21_28_port, QN => n_1675
               );
   REGISTERS_reg_21_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N157, next_state => N111, 
               clocked_on => CLK_port, Q => REGISTERS_21_27_port, QN => n_1676
               );
   REGISTERS_reg_21_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N157, next_state => N110, 
               clocked_on => CLK_port, Q => REGISTERS_21_26_port, QN => n_1677
               );
   REGISTERS_reg_21_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N157, next_state => N109, 
               clocked_on => CLK_port, Q => REGISTERS_21_25_port, QN => n_1678
               );
   REGISTERS_reg_21_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N157, next_state => N108, 
               clocked_on => CLK_port, Q => REGISTERS_21_24_port, QN => n_1679
               );
   REGISTERS_reg_21_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N157, next_state => N107, 
               clocked_on => CLK_port, Q => REGISTERS_21_23_port, QN => n_1680
               );
   REGISTERS_reg_21_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N157, next_state => N106, 
               clocked_on => CLK_port, Q => REGISTERS_21_22_port, QN => n_1681
               );
   REGISTERS_reg_21_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N157, next_state => N105, 
               clocked_on => CLK_port, Q => REGISTERS_21_21_port, QN => n_1682
               );
   REGISTERS_reg_21_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N157, next_state => N104, 
               clocked_on => CLK_port, Q => REGISTERS_21_20_port, QN => n_1683
               );
   REGISTERS_reg_21_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N157, next_state => N103, 
               clocked_on => CLK_port, Q => REGISTERS_21_19_port, QN => n_1684
               );
   REGISTERS_reg_21_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N157, next_state => N102, 
               clocked_on => CLK_port, Q => REGISTERS_21_18_port, QN => n_1685
               );
   REGISTERS_reg_21_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N157, next_state => N101, 
               clocked_on => CLK_port, Q => REGISTERS_21_17_port, QN => n_1686
               );
   REGISTERS_reg_21_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N157, next_state => N100, 
               clocked_on => CLK_port, Q => REGISTERS_21_16_port, QN => n_1687
               );
   REGISTERS_reg_21_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N157, next_state => N99, 
               clocked_on => CLK_port, Q => REGISTERS_21_15_port, QN => n_1688
               );
   REGISTERS_reg_21_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N157, next_state => N98, 
               clocked_on => CLK_port, Q => REGISTERS_21_14_port, QN => n_1689
               );
   REGISTERS_reg_21_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N157, next_state => N97, 
               clocked_on => CLK_port, Q => REGISTERS_21_13_port, QN => n_1690
               );
   REGISTERS_reg_21_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N157, next_state => N96, 
               clocked_on => CLK_port, Q => REGISTERS_21_12_port, QN => n_1691
               );
   REGISTERS_reg_21_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N157, next_state => N95, 
               clocked_on => CLK_port, Q => REGISTERS_21_11_port, QN => n_1692
               );
   REGISTERS_reg_21_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N157, next_state => N94, 
               clocked_on => CLK_port, Q => REGISTERS_21_10_port, QN => n_1693
               );
   REGISTERS_reg_21_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N157, next_state => N93, 
               clocked_on => CLK_port, Q => REGISTERS_21_9_port, QN => n_1694);
   REGISTERS_reg_21_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N157, next_state => N92, 
               clocked_on => CLK_port, Q => REGISTERS_21_8_port, QN => n_1695);
   REGISTERS_reg_21_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N157, next_state => N91, 
               clocked_on => CLK_port, Q => REGISTERS_21_7_port, QN => n_1696);
   REGISTERS_reg_21_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N157, next_state => N90, 
               clocked_on => CLK_port, Q => REGISTERS_21_6_port, QN => n_1697);
   REGISTERS_reg_21_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N157, next_state => N89, 
               clocked_on => CLK_port, Q => REGISTERS_21_5_port, QN => n_1698);
   REGISTERS_reg_21_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N157, next_state => N88, 
               clocked_on => CLK_port, Q => REGISTERS_21_4_port, QN => n_1699);
   REGISTERS_reg_21_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N157, next_state => N87, 
               clocked_on => CLK_port, Q => REGISTERS_21_3_port, QN => n_1700);
   REGISTERS_reg_21_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N157, next_state => N86, 
               clocked_on => CLK_port, Q => REGISTERS_21_2_port, QN => n_1701);
   REGISTERS_reg_21_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N157, next_state => N85, 
               clocked_on => CLK_port, Q => REGISTERS_21_1_port, QN => n_1702);
   REGISTERS_reg_21_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N157, next_state => N84, 
               clocked_on => CLK_port, Q => REGISTERS_21_0_port, QN => n_1703);
   REGISTERS_reg_22_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N156, next_state => N115, 
               clocked_on => CLK_port, Q => REGISTERS_22_31_port, QN => n_1704
               );
   REGISTERS_reg_22_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N156, next_state => N114, 
               clocked_on => CLK_port, Q => REGISTERS_22_30_port, QN => n_1705
               );
   REGISTERS_reg_22_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N156, next_state => N113, 
               clocked_on => CLK_port, Q => REGISTERS_22_29_port, QN => n_1706
               );
   REGISTERS_reg_22_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N156, next_state => N112, 
               clocked_on => CLK_port, Q => REGISTERS_22_28_port, QN => n_1707
               );
   REGISTERS_reg_22_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N156, next_state => N111, 
               clocked_on => CLK_port, Q => REGISTERS_22_27_port, QN => n_1708
               );
   REGISTERS_reg_22_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N156, next_state => N110, 
               clocked_on => CLK_port, Q => REGISTERS_22_26_port, QN => n_1709
               );
   REGISTERS_reg_22_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N156, next_state => N109, 
               clocked_on => CLK_port, Q => REGISTERS_22_25_port, QN => n_1710
               );
   REGISTERS_reg_22_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N156, next_state => N108, 
               clocked_on => CLK_port, Q => REGISTERS_22_24_port, QN => n_1711
               );
   REGISTERS_reg_22_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N156, next_state => N107, 
               clocked_on => CLK_port, Q => REGISTERS_22_23_port, QN => n_1712
               );
   REGISTERS_reg_22_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N156, next_state => N106, 
               clocked_on => CLK_port, Q => REGISTERS_22_22_port, QN => n_1713
               );
   REGISTERS_reg_22_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N156, next_state => N105, 
               clocked_on => CLK_port, Q => REGISTERS_22_21_port, QN => n_1714
               );
   REGISTERS_reg_22_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N156, next_state => N104, 
               clocked_on => CLK_port, Q => REGISTERS_22_20_port, QN => n_1715
               );
   REGISTERS_reg_22_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N156, next_state => N103, 
               clocked_on => CLK_port, Q => REGISTERS_22_19_port, QN => n_1716
               );
   REGISTERS_reg_22_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N156, next_state => N102, 
               clocked_on => CLK_port, Q => REGISTERS_22_18_port, QN => n_1717
               );
   REGISTERS_reg_22_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N156, next_state => N101, 
               clocked_on => CLK_port, Q => REGISTERS_22_17_port, QN => n_1718
               );
   REGISTERS_reg_22_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N156, next_state => N100, 
               clocked_on => CLK_port, Q => REGISTERS_22_16_port, QN => n_1719
               );
   REGISTERS_reg_22_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N156, next_state => N99, 
               clocked_on => CLK_port, Q => REGISTERS_22_15_port, QN => n_1720
               );
   REGISTERS_reg_22_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N156, next_state => N98, 
               clocked_on => CLK_port, Q => REGISTERS_22_14_port, QN => n_1721
               );
   REGISTERS_reg_22_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N156, next_state => N97, 
               clocked_on => CLK_port, Q => REGISTERS_22_13_port, QN => n_1722
               );
   REGISTERS_reg_22_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N156, next_state => N96, 
               clocked_on => CLK_port, Q => REGISTERS_22_12_port, QN => n_1723
               );
   REGISTERS_reg_22_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N156, next_state => N95, 
               clocked_on => CLK_port, Q => REGISTERS_22_11_port, QN => n_1724
               );
   REGISTERS_reg_22_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N156, next_state => N94, 
               clocked_on => CLK_port, Q => REGISTERS_22_10_port, QN => n_1725
               );
   REGISTERS_reg_22_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N156, next_state => N93, 
               clocked_on => CLK_port, Q => REGISTERS_22_9_port, QN => n_1726);
   REGISTERS_reg_22_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N156, next_state => N92, 
               clocked_on => CLK_port, Q => REGISTERS_22_8_port, QN => n_1727);
   REGISTERS_reg_22_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N156, next_state => N91, 
               clocked_on => CLK_port, Q => REGISTERS_22_7_port, QN => n_1728);
   REGISTERS_reg_22_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N156, next_state => N90, 
               clocked_on => CLK_port, Q => REGISTERS_22_6_port, QN => n_1729);
   REGISTERS_reg_22_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N156, next_state => N89, 
               clocked_on => CLK_port, Q => REGISTERS_22_5_port, QN => n_1730);
   REGISTERS_reg_22_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N156, next_state => N88, 
               clocked_on => CLK_port, Q => REGISTERS_22_4_port, QN => n_1731);
   REGISTERS_reg_22_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N156, next_state => N87, 
               clocked_on => CLK_port, Q => REGISTERS_22_3_port, QN => n_1732);
   REGISTERS_reg_22_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N156, next_state => N86, 
               clocked_on => CLK_port, Q => REGISTERS_22_2_port, QN => n_1733);
   REGISTERS_reg_22_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N156, next_state => N85, 
               clocked_on => CLK_port, Q => REGISTERS_22_1_port, QN => n_1734);
   REGISTERS_reg_22_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N156, next_state => N84, 
               clocked_on => CLK_port, Q => REGISTERS_22_0_port, QN => n_1735);
   REGISTERS_reg_23_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N155, next_state => N115, 
               clocked_on => CLK_port, Q => REGISTERS_23_31_port, QN => n_1736
               );
   REGISTERS_reg_23_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N155, next_state => N114, 
               clocked_on => CLK_port, Q => REGISTERS_23_30_port, QN => n_1737
               );
   REGISTERS_reg_23_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N155, next_state => N113, 
               clocked_on => CLK_port, Q => REGISTERS_23_29_port, QN => n_1738
               );
   REGISTERS_reg_23_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N155, next_state => N112, 
               clocked_on => CLK_port, Q => REGISTERS_23_28_port, QN => n_1739
               );
   REGISTERS_reg_23_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N155, next_state => N111, 
               clocked_on => CLK_port, Q => REGISTERS_23_27_port, QN => n_1740
               );
   REGISTERS_reg_23_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N155, next_state => N110, 
               clocked_on => CLK_port, Q => REGISTERS_23_26_port, QN => n_1741
               );
   REGISTERS_reg_23_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N155, next_state => N109, 
               clocked_on => CLK_port, Q => REGISTERS_23_25_port, QN => n_1742
               );
   REGISTERS_reg_23_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N155, next_state => N108, 
               clocked_on => CLK_port, Q => REGISTERS_23_24_port, QN => n_1743
               );
   REGISTERS_reg_23_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N155, next_state => N107, 
               clocked_on => CLK_port, Q => REGISTERS_23_23_port, QN => n_1744
               );
   REGISTERS_reg_23_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N155, next_state => N106, 
               clocked_on => CLK_port, Q => REGISTERS_23_22_port, QN => n_1745
               );
   REGISTERS_reg_23_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N155, next_state => N105, 
               clocked_on => CLK_port, Q => REGISTERS_23_21_port, QN => n_1746
               );
   REGISTERS_reg_23_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N155, next_state => N104, 
               clocked_on => CLK_port, Q => REGISTERS_23_20_port, QN => n_1747
               );
   REGISTERS_reg_23_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N155, next_state => N103, 
               clocked_on => CLK_port, Q => REGISTERS_23_19_port, QN => n_1748
               );
   REGISTERS_reg_23_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N155, next_state => N102, 
               clocked_on => CLK_port, Q => REGISTERS_23_18_port, QN => n_1749
               );
   REGISTERS_reg_23_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N155, next_state => N101, 
               clocked_on => CLK_port, Q => REGISTERS_23_17_port, QN => n_1750
               );
   REGISTERS_reg_23_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N155, next_state => N100, 
               clocked_on => CLK_port, Q => REGISTERS_23_16_port, QN => n_1751
               );
   REGISTERS_reg_23_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N155, next_state => N99, 
               clocked_on => CLK_port, Q => REGISTERS_23_15_port, QN => n_1752
               );
   REGISTERS_reg_23_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N155, next_state => N98, 
               clocked_on => CLK_port, Q => REGISTERS_23_14_port, QN => n_1753
               );
   REGISTERS_reg_23_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N155, next_state => N97, 
               clocked_on => CLK_port, Q => REGISTERS_23_13_port, QN => n_1754
               );
   REGISTERS_reg_23_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N155, next_state => N96, 
               clocked_on => CLK_port, Q => REGISTERS_23_12_port, QN => n_1755
               );
   REGISTERS_reg_23_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N155, next_state => N95, 
               clocked_on => CLK_port, Q => REGISTERS_23_11_port, QN => n_1756
               );
   REGISTERS_reg_23_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N155, next_state => N94, 
               clocked_on => CLK_port, Q => REGISTERS_23_10_port, QN => n_1757
               );
   REGISTERS_reg_23_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N155, next_state => N93, 
               clocked_on => CLK_port, Q => REGISTERS_23_9_port, QN => n_1758);
   REGISTERS_reg_23_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N155, next_state => N92, 
               clocked_on => CLK_port, Q => REGISTERS_23_8_port, QN => n_1759);
   REGISTERS_reg_23_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N155, next_state => N91, 
               clocked_on => CLK_port, Q => REGISTERS_23_7_port, QN => n_1760);
   REGISTERS_reg_23_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N155, next_state => N90, 
               clocked_on => CLK_port, Q => REGISTERS_23_6_port, QN => n_1761);
   REGISTERS_reg_23_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N155, next_state => N89, 
               clocked_on => CLK_port, Q => REGISTERS_23_5_port, QN => n_1762);
   REGISTERS_reg_23_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N155, next_state => N88, 
               clocked_on => CLK_port, Q => REGISTERS_23_4_port, QN => n_1763);
   REGISTERS_reg_23_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N155, next_state => N87, 
               clocked_on => CLK_port, Q => REGISTERS_23_3_port, QN => n_1764);
   REGISTERS_reg_23_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N155, next_state => N86, 
               clocked_on => CLK_port, Q => REGISTERS_23_2_port, QN => n_1765);
   REGISTERS_reg_23_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N155, next_state => N85, 
               clocked_on => CLK_port, Q => REGISTERS_23_1_port, QN => n_1766);
   REGISTERS_reg_23_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N155, next_state => N84, 
               clocked_on => CLK_port, Q => REGISTERS_23_0_port, QN => n_1767);
   REGISTERS_reg_24_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N154, next_state => N115, 
               clocked_on => CLK_port, Q => REGISTERS_24_31_port, QN => n_1768
               );
   REGISTERS_reg_24_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N154, next_state => N114, 
               clocked_on => CLK_port, Q => REGISTERS_24_30_port, QN => n_1769
               );
   REGISTERS_reg_24_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N154, next_state => N113, 
               clocked_on => CLK_port, Q => REGISTERS_24_29_port, QN => n_1770
               );
   REGISTERS_reg_24_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N154, next_state => N112, 
               clocked_on => CLK_port, Q => REGISTERS_24_28_port, QN => n_1771
               );
   REGISTERS_reg_24_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N154, next_state => N111, 
               clocked_on => CLK_port, Q => REGISTERS_24_27_port, QN => n_1772
               );
   REGISTERS_reg_24_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N154, next_state => N110, 
               clocked_on => CLK_port, Q => REGISTERS_24_26_port, QN => n_1773
               );
   REGISTERS_reg_24_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N154, next_state => N109, 
               clocked_on => CLK_port, Q => REGISTERS_24_25_port, QN => n_1774
               );
   REGISTERS_reg_24_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N154, next_state => N108, 
               clocked_on => CLK_port, Q => REGISTERS_24_24_port, QN => n_1775
               );
   REGISTERS_reg_24_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N154, next_state => N107, 
               clocked_on => CLK_port, Q => REGISTERS_24_23_port, QN => n_1776
               );
   REGISTERS_reg_24_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N154, next_state => N106, 
               clocked_on => CLK_port, Q => REGISTERS_24_22_port, QN => n_1777
               );
   REGISTERS_reg_24_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N154, next_state => N105, 
               clocked_on => CLK_port, Q => REGISTERS_24_21_port, QN => n_1778
               );
   REGISTERS_reg_24_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N154, next_state => N104, 
               clocked_on => CLK_port, Q => REGISTERS_24_20_port, QN => n_1779
               );
   REGISTERS_reg_24_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N154, next_state => N103, 
               clocked_on => CLK_port, Q => REGISTERS_24_19_port, QN => n_1780
               );
   REGISTERS_reg_24_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N154, next_state => N102, 
               clocked_on => CLK_port, Q => REGISTERS_24_18_port, QN => n_1781
               );
   REGISTERS_reg_24_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N154, next_state => N101, 
               clocked_on => CLK_port, Q => REGISTERS_24_17_port, QN => n_1782
               );
   REGISTERS_reg_24_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N154, next_state => N100, 
               clocked_on => CLK_port, Q => REGISTERS_24_16_port, QN => n_1783
               );
   REGISTERS_reg_24_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N154, next_state => N99, 
               clocked_on => CLK_port, Q => REGISTERS_24_15_port, QN => n_1784
               );
   REGISTERS_reg_24_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N154, next_state => N98, 
               clocked_on => CLK_port, Q => REGISTERS_24_14_port, QN => n_1785
               );
   REGISTERS_reg_24_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N154, next_state => N97, 
               clocked_on => CLK_port, Q => REGISTERS_24_13_port, QN => n_1786
               );
   REGISTERS_reg_24_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N154, next_state => N96, 
               clocked_on => CLK_port, Q => REGISTERS_24_12_port, QN => n_1787
               );
   REGISTERS_reg_24_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N154, next_state => N95, 
               clocked_on => CLK_port, Q => REGISTERS_24_11_port, QN => n_1788
               );
   REGISTERS_reg_24_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N154, next_state => N94, 
               clocked_on => CLK_port, Q => REGISTERS_24_10_port, QN => n_1789
               );
   REGISTERS_reg_24_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N154, next_state => N93, 
               clocked_on => CLK_port, Q => REGISTERS_24_9_port, QN => n_1790);
   REGISTERS_reg_24_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N154, next_state => N92, 
               clocked_on => CLK_port, Q => REGISTERS_24_8_port, QN => n_1791);
   REGISTERS_reg_24_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N154, next_state => N91, 
               clocked_on => CLK_port, Q => REGISTERS_24_7_port, QN => n_1792);
   REGISTERS_reg_24_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N154, next_state => N90, 
               clocked_on => CLK_port, Q => REGISTERS_24_6_port, QN => n_1793);
   REGISTERS_reg_24_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N154, next_state => N89, 
               clocked_on => CLK_port, Q => REGISTERS_24_5_port, QN => n_1794);
   REGISTERS_reg_24_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N154, next_state => N88, 
               clocked_on => CLK_port, Q => REGISTERS_24_4_port, QN => n_1795);
   REGISTERS_reg_24_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N154, next_state => N87, 
               clocked_on => CLK_port, Q => REGISTERS_24_3_port, QN => n_1796);
   REGISTERS_reg_24_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N154, next_state => N86, 
               clocked_on => CLK_port, Q => REGISTERS_24_2_port, QN => n_1797);
   REGISTERS_reg_24_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N154, next_state => N85, 
               clocked_on => CLK_port, Q => REGISTERS_24_1_port, QN => n_1798);
   REGISTERS_reg_24_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N154, next_state => N84, 
               clocked_on => CLK_port, Q => REGISTERS_24_0_port, QN => n_1799);
   REGISTERS_reg_25_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N153, next_state => N115, 
               clocked_on => CLK_port, Q => REGISTERS_25_31_port, QN => n_1800
               );
   REGISTERS_reg_25_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N153, next_state => N114, 
               clocked_on => CLK_port, Q => REGISTERS_25_30_port, QN => n_1801
               );
   REGISTERS_reg_25_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N153, next_state => N113, 
               clocked_on => CLK_port, Q => REGISTERS_25_29_port, QN => n_1802
               );
   REGISTERS_reg_25_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N153, next_state => N112, 
               clocked_on => CLK_port, Q => REGISTERS_25_28_port, QN => n_1803
               );
   REGISTERS_reg_25_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N153, next_state => N111, 
               clocked_on => CLK_port, Q => REGISTERS_25_27_port, QN => n_1804
               );
   REGISTERS_reg_25_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N153, next_state => N110, 
               clocked_on => CLK_port, Q => REGISTERS_25_26_port, QN => n_1805
               );
   REGISTERS_reg_25_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N153, next_state => N109, 
               clocked_on => CLK_port, Q => REGISTERS_25_25_port, QN => n_1806
               );
   REGISTERS_reg_25_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N153, next_state => N108, 
               clocked_on => CLK_port, Q => REGISTERS_25_24_port, QN => n_1807
               );
   REGISTERS_reg_25_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N153, next_state => N107, 
               clocked_on => CLK_port, Q => REGISTERS_25_23_port, QN => n_1808
               );
   REGISTERS_reg_25_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N153, next_state => N106, 
               clocked_on => CLK_port, Q => REGISTERS_25_22_port, QN => n_1809
               );
   REGISTERS_reg_25_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N153, next_state => N105, 
               clocked_on => CLK_port, Q => REGISTERS_25_21_port, QN => n_1810
               );
   REGISTERS_reg_25_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N153, next_state => N104, 
               clocked_on => CLK_port, Q => REGISTERS_25_20_port, QN => n_1811
               );
   REGISTERS_reg_25_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N153, next_state => N103, 
               clocked_on => CLK_port, Q => REGISTERS_25_19_port, QN => n_1812
               );
   REGISTERS_reg_25_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N153, next_state => N102, 
               clocked_on => CLK_port, Q => REGISTERS_25_18_port, QN => n_1813
               );
   REGISTERS_reg_25_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N153, next_state => N101, 
               clocked_on => CLK_port, Q => REGISTERS_25_17_port, QN => n_1814
               );
   REGISTERS_reg_25_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N153, next_state => N100, 
               clocked_on => CLK_port, Q => REGISTERS_25_16_port, QN => n_1815
               );
   REGISTERS_reg_25_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N153, next_state => N99, 
               clocked_on => CLK_port, Q => REGISTERS_25_15_port, QN => n_1816
               );
   REGISTERS_reg_25_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N153, next_state => N98, 
               clocked_on => CLK_port, Q => REGISTERS_25_14_port, QN => n_1817
               );
   REGISTERS_reg_25_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N153, next_state => N97, 
               clocked_on => CLK_port, Q => REGISTERS_25_13_port, QN => n_1818
               );
   REGISTERS_reg_25_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N153, next_state => N96, 
               clocked_on => CLK_port, Q => REGISTERS_25_12_port, QN => n_1819
               );
   REGISTERS_reg_25_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N153, next_state => N95, 
               clocked_on => CLK_port, Q => REGISTERS_25_11_port, QN => n_1820
               );
   REGISTERS_reg_25_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N153, next_state => N94, 
               clocked_on => CLK_port, Q => REGISTERS_25_10_port, QN => n_1821
               );
   REGISTERS_reg_25_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N153, next_state => N93, 
               clocked_on => CLK_port, Q => REGISTERS_25_9_port, QN => n_1822);
   REGISTERS_reg_25_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N153, next_state => N92, 
               clocked_on => CLK_port, Q => REGISTERS_25_8_port, QN => n_1823);
   REGISTERS_reg_25_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N153, next_state => N91, 
               clocked_on => CLK_port, Q => REGISTERS_25_7_port, QN => n_1824);
   REGISTERS_reg_25_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N153, next_state => N90, 
               clocked_on => CLK_port, Q => REGISTERS_25_6_port, QN => n_1825);
   REGISTERS_reg_25_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N153, next_state => N89, 
               clocked_on => CLK_port, Q => REGISTERS_25_5_port, QN => n_1826);
   REGISTERS_reg_25_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N153, next_state => N88, 
               clocked_on => CLK_port, Q => REGISTERS_25_4_port, QN => n_1827);
   REGISTERS_reg_25_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N153, next_state => N87, 
               clocked_on => CLK_port, Q => REGISTERS_25_3_port, QN => n_1828);
   REGISTERS_reg_25_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N153, next_state => N86, 
               clocked_on => CLK_port, Q => REGISTERS_25_2_port, QN => n_1829);
   REGISTERS_reg_25_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N153, next_state => N85, 
               clocked_on => CLK_port, Q => REGISTERS_25_1_port, QN => n_1830);
   REGISTERS_reg_25_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N153, next_state => N84, 
               clocked_on => CLK_port, Q => REGISTERS_25_0_port, QN => n_1831);
   REGISTERS_reg_26_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N152, next_state => N115, 
               clocked_on => CLK_port, Q => REGISTERS_26_31_port, QN => n_1832
               );
   REGISTERS_reg_26_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N152, next_state => N114, 
               clocked_on => CLK_port, Q => REGISTERS_26_30_port, QN => n_1833
               );
   REGISTERS_reg_26_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N152, next_state => N113, 
               clocked_on => CLK_port, Q => REGISTERS_26_29_port, QN => n_1834
               );
   REGISTERS_reg_26_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N152, next_state => N112, 
               clocked_on => CLK_port, Q => REGISTERS_26_28_port, QN => n_1835
               );
   REGISTERS_reg_26_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N152, next_state => N111, 
               clocked_on => CLK_port, Q => REGISTERS_26_27_port, QN => n_1836
               );
   REGISTERS_reg_26_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N152, next_state => N110, 
               clocked_on => CLK_port, Q => REGISTERS_26_26_port, QN => n_1837
               );
   REGISTERS_reg_26_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N152, next_state => N109, 
               clocked_on => CLK_port, Q => REGISTERS_26_25_port, QN => n_1838
               );
   REGISTERS_reg_26_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N152, next_state => N108, 
               clocked_on => CLK_port, Q => REGISTERS_26_24_port, QN => n_1839
               );
   REGISTERS_reg_26_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N152, next_state => N107, 
               clocked_on => CLK_port, Q => REGISTERS_26_23_port, QN => n_1840
               );
   REGISTERS_reg_26_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N152, next_state => N106, 
               clocked_on => CLK_port, Q => REGISTERS_26_22_port, QN => n_1841
               );
   REGISTERS_reg_26_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N152, next_state => N105, 
               clocked_on => CLK_port, Q => REGISTERS_26_21_port, QN => n_1842
               );
   REGISTERS_reg_26_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N152, next_state => N104, 
               clocked_on => CLK_port, Q => REGISTERS_26_20_port, QN => n_1843
               );
   REGISTERS_reg_26_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N152, next_state => N103, 
               clocked_on => CLK_port, Q => REGISTERS_26_19_port, QN => n_1844
               );
   REGISTERS_reg_26_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N152, next_state => N102, 
               clocked_on => CLK_port, Q => REGISTERS_26_18_port, QN => n_1845
               );
   REGISTERS_reg_26_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N152, next_state => N101, 
               clocked_on => CLK_port, Q => REGISTERS_26_17_port, QN => n_1846
               );
   REGISTERS_reg_26_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N152, next_state => N100, 
               clocked_on => CLK_port, Q => REGISTERS_26_16_port, QN => n_1847
               );
   REGISTERS_reg_26_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N152, next_state => N99, 
               clocked_on => CLK_port, Q => REGISTERS_26_15_port, QN => n_1848
               );
   REGISTERS_reg_26_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N152, next_state => N98, 
               clocked_on => CLK_port, Q => REGISTERS_26_14_port, QN => n_1849
               );
   REGISTERS_reg_26_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N152, next_state => N97, 
               clocked_on => CLK_port, Q => REGISTERS_26_13_port, QN => n_1850
               );
   REGISTERS_reg_26_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N152, next_state => N96, 
               clocked_on => CLK_port, Q => REGISTERS_26_12_port, QN => n_1851
               );
   REGISTERS_reg_26_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N152, next_state => N95, 
               clocked_on => CLK_port, Q => REGISTERS_26_11_port, QN => n_1852
               );
   REGISTERS_reg_26_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N152, next_state => N94, 
               clocked_on => CLK_port, Q => REGISTERS_26_10_port, QN => n_1853
               );
   REGISTERS_reg_26_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N152, next_state => N93, 
               clocked_on => CLK_port, Q => REGISTERS_26_9_port, QN => n_1854);
   REGISTERS_reg_26_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N152, next_state => N92, 
               clocked_on => CLK_port, Q => REGISTERS_26_8_port, QN => n_1855);
   REGISTERS_reg_26_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N152, next_state => N91, 
               clocked_on => CLK_port, Q => REGISTERS_26_7_port, QN => n_1856);
   REGISTERS_reg_26_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N152, next_state => N90, 
               clocked_on => CLK_port, Q => REGISTERS_26_6_port, QN => n_1857);
   REGISTERS_reg_26_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N152, next_state => N89, 
               clocked_on => CLK_port, Q => REGISTERS_26_5_port, QN => n_1858);
   REGISTERS_reg_26_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N152, next_state => N88, 
               clocked_on => CLK_port, Q => REGISTERS_26_4_port, QN => n_1859);
   REGISTERS_reg_26_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N152, next_state => N87, 
               clocked_on => CLK_port, Q => REGISTERS_26_3_port, QN => n_1860);
   REGISTERS_reg_26_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N152, next_state => N86, 
               clocked_on => CLK_port, Q => REGISTERS_26_2_port, QN => n_1861);
   REGISTERS_reg_26_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N152, next_state => N85, 
               clocked_on => CLK_port, Q => REGISTERS_26_1_port, QN => n_1862);
   REGISTERS_reg_26_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N152, next_state => N84, 
               clocked_on => CLK_port, Q => REGISTERS_26_0_port, QN => n_1863);
   REGISTERS_reg_27_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N151, next_state => N115, 
               clocked_on => CLK_port, Q => REGISTERS_27_31_port, QN => n_1864
               );
   REGISTERS_reg_27_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N151, next_state => N114, 
               clocked_on => CLK_port, Q => REGISTERS_27_30_port, QN => n_1865
               );
   REGISTERS_reg_27_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N151, next_state => N113, 
               clocked_on => CLK_port, Q => REGISTERS_27_29_port, QN => n_1866
               );
   REGISTERS_reg_27_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N151, next_state => N112, 
               clocked_on => CLK_port, Q => REGISTERS_27_28_port, QN => n_1867
               );
   REGISTERS_reg_27_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N151, next_state => N111, 
               clocked_on => CLK_port, Q => REGISTERS_27_27_port, QN => n_1868
               );
   REGISTERS_reg_27_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N151, next_state => N110, 
               clocked_on => CLK_port, Q => REGISTERS_27_26_port, QN => n_1869
               );
   REGISTERS_reg_27_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N151, next_state => N109, 
               clocked_on => CLK_port, Q => REGISTERS_27_25_port, QN => n_1870
               );
   REGISTERS_reg_27_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N151, next_state => N108, 
               clocked_on => CLK_port, Q => REGISTERS_27_24_port, QN => n_1871
               );
   REGISTERS_reg_27_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N151, next_state => N107, 
               clocked_on => CLK_port, Q => REGISTERS_27_23_port, QN => n_1872
               );
   REGISTERS_reg_27_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N151, next_state => N106, 
               clocked_on => CLK_port, Q => REGISTERS_27_22_port, QN => n_1873
               );
   REGISTERS_reg_27_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N151, next_state => N105, 
               clocked_on => CLK_port, Q => REGISTERS_27_21_port, QN => n_1874
               );
   REGISTERS_reg_27_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N151, next_state => N104, 
               clocked_on => CLK_port, Q => REGISTERS_27_20_port, QN => n_1875
               );
   REGISTERS_reg_27_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N151, next_state => N103, 
               clocked_on => CLK_port, Q => REGISTERS_27_19_port, QN => n_1876
               );
   REGISTERS_reg_27_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N151, next_state => N102, 
               clocked_on => CLK_port, Q => REGISTERS_27_18_port, QN => n_1877
               );
   REGISTERS_reg_27_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N151, next_state => N101, 
               clocked_on => CLK_port, Q => REGISTERS_27_17_port, QN => n_1878
               );
   REGISTERS_reg_27_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N151, next_state => N100, 
               clocked_on => CLK_port, Q => REGISTERS_27_16_port, QN => n_1879
               );
   REGISTERS_reg_27_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N151, next_state => N99, 
               clocked_on => CLK_port, Q => REGISTERS_27_15_port, QN => n_1880
               );
   REGISTERS_reg_27_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N151, next_state => N98, 
               clocked_on => CLK_port, Q => REGISTERS_27_14_port, QN => n_1881
               );
   REGISTERS_reg_27_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N151, next_state => N97, 
               clocked_on => CLK_port, Q => REGISTERS_27_13_port, QN => n_1882
               );
   REGISTERS_reg_27_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N151, next_state => N96, 
               clocked_on => CLK_port, Q => REGISTERS_27_12_port, QN => n_1883
               );
   REGISTERS_reg_27_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N151, next_state => N95, 
               clocked_on => CLK_port, Q => REGISTERS_27_11_port, QN => n_1884
               );
   REGISTERS_reg_27_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N151, next_state => N94, 
               clocked_on => CLK_port, Q => REGISTERS_27_10_port, QN => n_1885
               );
   REGISTERS_reg_27_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N151, next_state => N93, 
               clocked_on => CLK_port, Q => REGISTERS_27_9_port, QN => n_1886);
   REGISTERS_reg_27_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N151, next_state => N92, 
               clocked_on => CLK_port, Q => REGISTERS_27_8_port, QN => n_1887);
   REGISTERS_reg_27_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N151, next_state => N91, 
               clocked_on => CLK_port, Q => REGISTERS_27_7_port, QN => n_1888);
   REGISTERS_reg_27_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N151, next_state => N90, 
               clocked_on => CLK_port, Q => REGISTERS_27_6_port, QN => n_1889);
   REGISTERS_reg_27_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N151, next_state => N89, 
               clocked_on => CLK_port, Q => REGISTERS_27_5_port, QN => n_1890);
   REGISTERS_reg_27_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N151, next_state => N88, 
               clocked_on => CLK_port, Q => REGISTERS_27_4_port, QN => n_1891);
   REGISTERS_reg_27_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N151, next_state => N87, 
               clocked_on => CLK_port, Q => REGISTERS_27_3_port, QN => n_1892);
   REGISTERS_reg_27_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N151, next_state => N86, 
               clocked_on => CLK_port, Q => REGISTERS_27_2_port, QN => n_1893);
   REGISTERS_reg_27_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N151, next_state => N85, 
               clocked_on => CLK_port, Q => REGISTERS_27_1_port, QN => n_1894);
   REGISTERS_reg_27_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N151, next_state => N84, 
               clocked_on => CLK_port, Q => REGISTERS_27_0_port, QN => n_1895);
   REGISTERS_reg_28_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N150, next_state => N115, 
               clocked_on => CLK_port, Q => REGISTERS_28_31_port, QN => n_1896
               );
   REGISTERS_reg_28_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N150, next_state => N114, 
               clocked_on => CLK_port, Q => REGISTERS_28_30_port, QN => n_1897
               );
   REGISTERS_reg_28_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N150, next_state => N113, 
               clocked_on => CLK_port, Q => REGISTERS_28_29_port, QN => n_1898
               );
   REGISTERS_reg_28_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N150, next_state => N112, 
               clocked_on => CLK_port, Q => REGISTERS_28_28_port, QN => n_1899
               );
   REGISTERS_reg_28_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N150, next_state => N111, 
               clocked_on => CLK_port, Q => REGISTERS_28_27_port, QN => n_1900
               );
   REGISTERS_reg_28_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N150, next_state => N110, 
               clocked_on => CLK_port, Q => REGISTERS_28_26_port, QN => n_1901
               );
   REGISTERS_reg_28_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N150, next_state => N109, 
               clocked_on => CLK_port, Q => REGISTERS_28_25_port, QN => n_1902
               );
   REGISTERS_reg_28_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N150, next_state => N108, 
               clocked_on => CLK_port, Q => REGISTERS_28_24_port, QN => n_1903
               );
   REGISTERS_reg_28_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N150, next_state => N107, 
               clocked_on => CLK_port, Q => REGISTERS_28_23_port, QN => n_1904
               );
   REGISTERS_reg_28_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N150, next_state => N106, 
               clocked_on => CLK_port, Q => REGISTERS_28_22_port, QN => n_1905
               );
   REGISTERS_reg_28_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N150, next_state => N105, 
               clocked_on => CLK_port, Q => REGISTERS_28_21_port, QN => n_1906
               );
   REGISTERS_reg_28_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N150, next_state => N104, 
               clocked_on => CLK_port, Q => REGISTERS_28_20_port, QN => n_1907
               );
   REGISTERS_reg_28_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N150, next_state => N103, 
               clocked_on => CLK_port, Q => REGISTERS_28_19_port, QN => n_1908
               );
   REGISTERS_reg_28_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N150, next_state => N102, 
               clocked_on => CLK_port, Q => REGISTERS_28_18_port, QN => n_1909
               );
   REGISTERS_reg_28_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N150, next_state => N101, 
               clocked_on => CLK_port, Q => REGISTERS_28_17_port, QN => n_1910
               );
   REGISTERS_reg_28_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N150, next_state => N100, 
               clocked_on => CLK_port, Q => REGISTERS_28_16_port, QN => n_1911
               );
   REGISTERS_reg_28_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N150, next_state => N99, 
               clocked_on => CLK_port, Q => REGISTERS_28_15_port, QN => n_1912
               );
   REGISTERS_reg_28_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N150, next_state => N98, 
               clocked_on => CLK_port, Q => REGISTERS_28_14_port, QN => n_1913
               );
   REGISTERS_reg_28_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N150, next_state => N97, 
               clocked_on => CLK_port, Q => REGISTERS_28_13_port, QN => n_1914
               );
   REGISTERS_reg_28_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N150, next_state => N96, 
               clocked_on => CLK_port, Q => REGISTERS_28_12_port, QN => n_1915
               );
   REGISTERS_reg_28_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N150, next_state => N95, 
               clocked_on => CLK_port, Q => REGISTERS_28_11_port, QN => n_1916
               );
   REGISTERS_reg_28_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N150, next_state => N94, 
               clocked_on => CLK_port, Q => REGISTERS_28_10_port, QN => n_1917
               );
   REGISTERS_reg_28_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N150, next_state => N93, 
               clocked_on => CLK_port, Q => REGISTERS_28_9_port, QN => n_1918);
   REGISTERS_reg_28_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N150, next_state => N92, 
               clocked_on => CLK_port, Q => REGISTERS_28_8_port, QN => n_1919);
   REGISTERS_reg_28_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N150, next_state => N91, 
               clocked_on => CLK_port, Q => REGISTERS_28_7_port, QN => n_1920);
   REGISTERS_reg_28_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N150, next_state => N90, 
               clocked_on => CLK_port, Q => REGISTERS_28_6_port, QN => n_1921);
   REGISTERS_reg_28_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N150, next_state => N89, 
               clocked_on => CLK_port, Q => REGISTERS_28_5_port, QN => n_1922);
   REGISTERS_reg_28_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N150, next_state => N88, 
               clocked_on => CLK_port, Q => REGISTERS_28_4_port, QN => n_1923);
   REGISTERS_reg_28_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N150, next_state => N87, 
               clocked_on => CLK_port, Q => REGISTERS_28_3_port, QN => n_1924);
   REGISTERS_reg_28_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N150, next_state => N86, 
               clocked_on => CLK_port, Q => REGISTERS_28_2_port, QN => n_1925);
   REGISTERS_reg_28_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N150, next_state => N85, 
               clocked_on => CLK_port, Q => REGISTERS_28_1_port, QN => n_1926);
   REGISTERS_reg_28_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N150, next_state => N84, 
               clocked_on => CLK_port, Q => REGISTERS_28_0_port, QN => n_1927);
   REGISTERS_reg_29_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N149, next_state => N115, 
               clocked_on => CLK_port, Q => REGISTERS_29_31_port, QN => n_1928
               );
   REGISTERS_reg_29_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N149, next_state => N114, 
               clocked_on => CLK_port, Q => REGISTERS_29_30_port, QN => n_1929
               );
   REGISTERS_reg_29_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N149, next_state => N113, 
               clocked_on => CLK_port, Q => REGISTERS_29_29_port, QN => n_1930
               );
   REGISTERS_reg_29_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N149, next_state => N112, 
               clocked_on => CLK_port, Q => REGISTERS_29_28_port, QN => n_1931
               );
   REGISTERS_reg_29_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N149, next_state => N111, 
               clocked_on => CLK_port, Q => REGISTERS_29_27_port, QN => n_1932
               );
   REGISTERS_reg_29_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N149, next_state => N110, 
               clocked_on => CLK_port, Q => REGISTERS_29_26_port, QN => n_1933
               );
   REGISTERS_reg_29_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N149, next_state => N109, 
               clocked_on => CLK_port, Q => REGISTERS_29_25_port, QN => n_1934
               );
   REGISTERS_reg_29_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N149, next_state => N108, 
               clocked_on => CLK_port, Q => REGISTERS_29_24_port, QN => n_1935
               );
   REGISTERS_reg_29_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N149, next_state => N107, 
               clocked_on => CLK_port, Q => REGISTERS_29_23_port, QN => n_1936
               );
   REGISTERS_reg_29_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N149, next_state => N106, 
               clocked_on => CLK_port, Q => REGISTERS_29_22_port, QN => n_1937
               );
   REGISTERS_reg_29_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N149, next_state => N105, 
               clocked_on => CLK_port, Q => REGISTERS_29_21_port, QN => n_1938
               );
   REGISTERS_reg_29_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N149, next_state => N104, 
               clocked_on => CLK_port, Q => REGISTERS_29_20_port, QN => n_1939
               );
   REGISTERS_reg_29_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N149, next_state => N103, 
               clocked_on => CLK_port, Q => REGISTERS_29_19_port, QN => n_1940
               );
   REGISTERS_reg_29_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N149, next_state => N102, 
               clocked_on => CLK_port, Q => REGISTERS_29_18_port, QN => n_1941
               );
   REGISTERS_reg_29_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N149, next_state => N101, 
               clocked_on => CLK_port, Q => REGISTERS_29_17_port, QN => n_1942
               );
   REGISTERS_reg_29_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N149, next_state => N100, 
               clocked_on => CLK_port, Q => REGISTERS_29_16_port, QN => n_1943
               );
   REGISTERS_reg_29_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N149, next_state => N99, 
               clocked_on => CLK_port, Q => REGISTERS_29_15_port, QN => n_1944
               );
   REGISTERS_reg_29_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N149, next_state => N98, 
               clocked_on => CLK_port, Q => REGISTERS_29_14_port, QN => n_1945
               );
   REGISTERS_reg_29_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N149, next_state => N97, 
               clocked_on => CLK_port, Q => REGISTERS_29_13_port, QN => n_1946
               );
   REGISTERS_reg_29_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N149, next_state => N96, 
               clocked_on => CLK_port, Q => REGISTERS_29_12_port, QN => n_1947
               );
   REGISTERS_reg_29_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N149, next_state => N95, 
               clocked_on => CLK_port, Q => REGISTERS_29_11_port, QN => n_1948
               );
   REGISTERS_reg_29_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N149, next_state => N94, 
               clocked_on => CLK_port, Q => REGISTERS_29_10_port, QN => n_1949
               );
   REGISTERS_reg_29_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N149, next_state => N93, 
               clocked_on => CLK_port, Q => REGISTERS_29_9_port, QN => n_1950);
   REGISTERS_reg_29_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N149, next_state => N92, 
               clocked_on => CLK_port, Q => REGISTERS_29_8_port, QN => n_1951);
   REGISTERS_reg_29_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N149, next_state => N91, 
               clocked_on => CLK_port, Q => REGISTERS_29_7_port, QN => n_1952);
   REGISTERS_reg_29_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N149, next_state => N90, 
               clocked_on => CLK_port, Q => REGISTERS_29_6_port, QN => n_1953);
   REGISTERS_reg_29_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N149, next_state => N89, 
               clocked_on => CLK_port, Q => REGISTERS_29_5_port, QN => n_1954);
   REGISTERS_reg_29_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N149, next_state => N88, 
               clocked_on => CLK_port, Q => REGISTERS_29_4_port, QN => n_1955);
   REGISTERS_reg_29_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N149, next_state => N87, 
               clocked_on => CLK_port, Q => REGISTERS_29_3_port, QN => n_1956);
   REGISTERS_reg_29_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N149, next_state => N86, 
               clocked_on => CLK_port, Q => REGISTERS_29_2_port, QN => n_1957);
   REGISTERS_reg_29_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N149, next_state => N85, 
               clocked_on => CLK_port, Q => REGISTERS_29_1_port, QN => n_1958);
   REGISTERS_reg_29_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N149, next_state => N84, 
               clocked_on => CLK_port, Q => REGISTERS_29_0_port, QN => n_1959);
   REGISTERS_reg_30_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N148, next_state => N115, 
               clocked_on => CLK_port, Q => REGISTERS_30_31_port, QN => n_1960
               );
   REGISTERS_reg_30_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N148, next_state => N114, 
               clocked_on => CLK_port, Q => REGISTERS_30_30_port, QN => n_1961
               );
   REGISTERS_reg_30_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N148, next_state => N113, 
               clocked_on => CLK_port, Q => REGISTERS_30_29_port, QN => n_1962
               );
   REGISTERS_reg_30_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N148, next_state => N112, 
               clocked_on => CLK_port, Q => REGISTERS_30_28_port, QN => n_1963
               );
   REGISTERS_reg_30_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N148, next_state => N111, 
               clocked_on => CLK_port, Q => REGISTERS_30_27_port, QN => n_1964
               );
   REGISTERS_reg_30_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N148, next_state => N110, 
               clocked_on => CLK_port, Q => REGISTERS_30_26_port, QN => n_1965
               );
   REGISTERS_reg_30_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N148, next_state => N109, 
               clocked_on => CLK_port, Q => REGISTERS_30_25_port, QN => n_1966
               );
   REGISTERS_reg_30_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N148, next_state => N108, 
               clocked_on => CLK_port, Q => REGISTERS_30_24_port, QN => n_1967
               );
   REGISTERS_reg_30_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N148, next_state => N107, 
               clocked_on => CLK_port, Q => REGISTERS_30_23_port, QN => n_1968
               );
   REGISTERS_reg_30_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N148, next_state => N106, 
               clocked_on => CLK_port, Q => REGISTERS_30_22_port, QN => n_1969
               );
   REGISTERS_reg_30_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N148, next_state => N105, 
               clocked_on => CLK_port, Q => REGISTERS_30_21_port, QN => n_1970
               );
   REGISTERS_reg_30_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N148, next_state => N104, 
               clocked_on => CLK_port, Q => REGISTERS_30_20_port, QN => n_1971
               );
   REGISTERS_reg_30_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N148, next_state => N103, 
               clocked_on => CLK_port, Q => REGISTERS_30_19_port, QN => n_1972
               );
   REGISTERS_reg_30_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N148, next_state => N102, 
               clocked_on => CLK_port, Q => REGISTERS_30_18_port, QN => n_1973
               );
   REGISTERS_reg_30_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N148, next_state => N101, 
               clocked_on => CLK_port, Q => REGISTERS_30_17_port, QN => n_1974
               );
   REGISTERS_reg_30_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N148, next_state => N100, 
               clocked_on => CLK_port, Q => REGISTERS_30_16_port, QN => n_1975
               );
   REGISTERS_reg_30_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N148, next_state => N99, 
               clocked_on => CLK_port, Q => REGISTERS_30_15_port, QN => n_1976
               );
   REGISTERS_reg_30_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N148, next_state => N98, 
               clocked_on => CLK_port, Q => REGISTERS_30_14_port, QN => n_1977
               );
   REGISTERS_reg_30_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N148, next_state => N97, 
               clocked_on => CLK_port, Q => REGISTERS_30_13_port, QN => n_1978
               );
   REGISTERS_reg_30_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N148, next_state => N96, 
               clocked_on => CLK_port, Q => REGISTERS_30_12_port, QN => n_1979
               );
   REGISTERS_reg_30_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N148, next_state => N95, 
               clocked_on => CLK_port, Q => REGISTERS_30_11_port, QN => n_1980
               );
   REGISTERS_reg_30_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N148, next_state => N94, 
               clocked_on => CLK_port, Q => REGISTERS_30_10_port, QN => n_1981
               );
   REGISTERS_reg_30_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N148, next_state => N93, 
               clocked_on => CLK_port, Q => REGISTERS_30_9_port, QN => n_1982);
   REGISTERS_reg_30_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N148, next_state => N92, 
               clocked_on => CLK_port, Q => REGISTERS_30_8_port, QN => n_1983);
   REGISTERS_reg_30_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N148, next_state => N91, 
               clocked_on => CLK_port, Q => REGISTERS_30_7_port, QN => n_1984);
   REGISTERS_reg_30_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N148, next_state => N90, 
               clocked_on => CLK_port, Q => REGISTERS_30_6_port, QN => n_1985);
   REGISTERS_reg_30_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N148, next_state => N89, 
               clocked_on => CLK_port, Q => REGISTERS_30_5_port, QN => n_1986);
   REGISTERS_reg_30_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N148, next_state => N88, 
               clocked_on => CLK_port, Q => REGISTERS_30_4_port, QN => n_1987);
   REGISTERS_reg_30_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N148, next_state => N87, 
               clocked_on => CLK_port, Q => REGISTERS_30_3_port, QN => n_1988);
   REGISTERS_reg_30_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N148, next_state => N86, 
               clocked_on => CLK_port, Q => REGISTERS_30_2_port, QN => n_1989);
   REGISTERS_reg_30_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N148, next_state => N85, 
               clocked_on => CLK_port, Q => REGISTERS_30_1_port, QN => n_1990);
   REGISTERS_reg_30_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N148, next_state => N84, 
               clocked_on => CLK_port, Q => REGISTERS_30_0_port, QN => n_1991);
   REGISTERS_reg_31_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N147, next_state => N115, 
               clocked_on => CLK_port, Q => REGISTERS_31_31_port, QN => n_1992
               );
   REGISTERS_reg_31_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N147, next_state => N114, 
               clocked_on => CLK_port, Q => REGISTERS_31_30_port, QN => n_1993
               );
   REGISTERS_reg_31_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N147, next_state => N113, 
               clocked_on => CLK_port, Q => REGISTERS_31_29_port, QN => n_1994
               );
   REGISTERS_reg_31_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N147, next_state => N112, 
               clocked_on => CLK_port, Q => REGISTERS_31_28_port, QN => n_1995
               );
   REGISTERS_reg_31_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N147, next_state => N111, 
               clocked_on => CLK_port, Q => REGISTERS_31_27_port, QN => n_1996
               );
   REGISTERS_reg_31_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N147, next_state => N110, 
               clocked_on => CLK_port, Q => REGISTERS_31_26_port, QN => n_1997
               );
   REGISTERS_reg_31_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N147, next_state => N109, 
               clocked_on => CLK_port, Q => REGISTERS_31_25_port, QN => n_1998
               );
   REGISTERS_reg_31_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N147, next_state => N108, 
               clocked_on => CLK_port, Q => REGISTERS_31_24_port, QN => n_1999
               );
   REGISTERS_reg_31_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N147, next_state => N107, 
               clocked_on => CLK_port, Q => REGISTERS_31_23_port, QN => n_2000
               );
   REGISTERS_reg_31_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N147, next_state => N106, 
               clocked_on => CLK_port, Q => REGISTERS_31_22_port, QN => n_2001
               );
   REGISTERS_reg_31_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N147, next_state => N105, 
               clocked_on => CLK_port, Q => REGISTERS_31_21_port, QN => n_2002
               );
   REGISTERS_reg_31_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N147, next_state => N104, 
               clocked_on => CLK_port, Q => REGISTERS_31_20_port, QN => n_2003
               );
   REGISTERS_reg_31_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N147, next_state => N103, 
               clocked_on => CLK_port, Q => REGISTERS_31_19_port, QN => n_2004
               );
   REGISTERS_reg_31_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N147, next_state => N102, 
               clocked_on => CLK_port, Q => REGISTERS_31_18_port, QN => n_2005
               );
   REGISTERS_reg_31_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N147, next_state => N101, 
               clocked_on => CLK_port, Q => REGISTERS_31_17_port, QN => n_2006
               );
   REGISTERS_reg_31_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N147, next_state => N100, 
               clocked_on => CLK_port, Q => REGISTERS_31_16_port, QN => n_2007
               );
   REGISTERS_reg_31_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N147, next_state => N99, 
               clocked_on => CLK_port, Q => REGISTERS_31_15_port, QN => n_2008
               );
   REGISTERS_reg_31_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N147, next_state => N98, 
               clocked_on => CLK_port, Q => REGISTERS_31_14_port, QN => n_2009
               );
   REGISTERS_reg_31_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N147, next_state => N97, 
               clocked_on => CLK_port, Q => REGISTERS_31_13_port, QN => n_2010
               );
   REGISTERS_reg_31_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N147, next_state => N96, 
               clocked_on => CLK_port, Q => REGISTERS_31_12_port, QN => n_2011
               );
   REGISTERS_reg_31_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N147, next_state => N95, 
               clocked_on => CLK_port, Q => REGISTERS_31_11_port, QN => n_2012
               );
   REGISTERS_reg_31_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N147, next_state => N94, 
               clocked_on => CLK_port, Q => REGISTERS_31_10_port, QN => n_2013
               );
   REGISTERS_reg_31_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N147, next_state => N93, 
               clocked_on => CLK_port, Q => REGISTERS_31_9_port, QN => n_2014);
   REGISTERS_reg_31_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N147, next_state => N92, 
               clocked_on => CLK_port, Q => REGISTERS_31_8_port, QN => n_2015);
   REGISTERS_reg_31_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N147, next_state => N91, 
               clocked_on => CLK_port, Q => REGISTERS_31_7_port, QN => n_2016);
   REGISTERS_reg_31_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N147, next_state => N90, 
               clocked_on => CLK_port, Q => REGISTERS_31_6_port, QN => n_2017);
   REGISTERS_reg_31_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N147, next_state => N89, 
               clocked_on => CLK_port, Q => REGISTERS_31_5_port, QN => n_2018);
   REGISTERS_reg_31_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N147, next_state => N88, 
               clocked_on => CLK_port, Q => REGISTERS_31_4_port, QN => n_2019);
   REGISTERS_reg_31_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N147, next_state => N87, 
               clocked_on => CLK_port, Q => REGISTERS_31_3_port, QN => n_2020);
   REGISTERS_reg_31_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N147, next_state => N86, 
               clocked_on => CLK_port, Q => REGISTERS_31_2_port, QN => n_2021);
   REGISTERS_reg_31_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N147, next_state => N85, 
               clocked_on => CLK_port, Q => REGISTERS_31_1_port, QN => n_2022);
   REGISTERS_reg_31_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N147, next_state => N84, 
               clocked_on => CLK_port, Q => REGISTERS_31_0_port, QN => n_2023);
   REGISTERS_reg_32_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N146, next_state => N115, 
               clocked_on => CLK_port, Q => REGISTERS_32_31_port, QN => n_2024
               );
   REGISTERS_reg_32_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N146, next_state => N114, 
               clocked_on => CLK_port, Q => REGISTERS_32_30_port, QN => n_2025
               );
   REGISTERS_reg_32_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N146, next_state => N113, 
               clocked_on => CLK_port, Q => REGISTERS_32_29_port, QN => n_2026
               );
   REGISTERS_reg_32_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N146, next_state => N112, 
               clocked_on => CLK_port, Q => REGISTERS_32_28_port, QN => n_2027
               );
   REGISTERS_reg_32_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N146, next_state => N111, 
               clocked_on => CLK_port, Q => REGISTERS_32_27_port, QN => n_2028
               );
   REGISTERS_reg_32_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N146, next_state => N110, 
               clocked_on => CLK_port, Q => REGISTERS_32_26_port, QN => n_2029
               );
   REGISTERS_reg_32_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N146, next_state => N109, 
               clocked_on => CLK_port, Q => REGISTERS_32_25_port, QN => n_2030
               );
   REGISTERS_reg_32_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N146, next_state => N108, 
               clocked_on => CLK_port, Q => REGISTERS_32_24_port, QN => n_2031
               );
   REGISTERS_reg_32_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N146, next_state => N107, 
               clocked_on => CLK_port, Q => REGISTERS_32_23_port, QN => n_2032
               );
   REGISTERS_reg_32_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N146, next_state => N106, 
               clocked_on => CLK_port, Q => REGISTERS_32_22_port, QN => n_2033
               );
   REGISTERS_reg_32_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N146, next_state => N105, 
               clocked_on => CLK_port, Q => REGISTERS_32_21_port, QN => n_2034
               );
   REGISTERS_reg_32_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N146, next_state => N104, 
               clocked_on => CLK_port, Q => REGISTERS_32_20_port, QN => n_2035
               );
   REGISTERS_reg_32_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N146, next_state => N103, 
               clocked_on => CLK_port, Q => REGISTERS_32_19_port, QN => n_2036
               );
   REGISTERS_reg_32_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N146, next_state => N102, 
               clocked_on => CLK_port, Q => REGISTERS_32_18_port, QN => n_2037
               );
   REGISTERS_reg_32_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N146, next_state => N101, 
               clocked_on => CLK_port, Q => REGISTERS_32_17_port, QN => n_2038
               );
   REGISTERS_reg_32_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N146, next_state => N100, 
               clocked_on => CLK_port, Q => REGISTERS_32_16_port, QN => n_2039
               );
   REGISTERS_reg_32_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N146, next_state => N99, 
               clocked_on => CLK_port, Q => REGISTERS_32_15_port, QN => n_2040
               );
   REGISTERS_reg_32_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N146, next_state => N98, 
               clocked_on => CLK_port, Q => REGISTERS_32_14_port, QN => n_2041
               );
   REGISTERS_reg_32_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N146, next_state => N97, 
               clocked_on => CLK_port, Q => REGISTERS_32_13_port, QN => n_2042
               );
   REGISTERS_reg_32_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N146, next_state => N96, 
               clocked_on => CLK_port, Q => REGISTERS_32_12_port, QN => n_2043
               );
   REGISTERS_reg_32_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N146, next_state => N95, 
               clocked_on => CLK_port, Q => REGISTERS_32_11_port, QN => n_2044
               );
   REGISTERS_reg_32_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N146, next_state => N94, 
               clocked_on => CLK_port, Q => REGISTERS_32_10_port, QN => n_2045
               );
   REGISTERS_reg_32_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N146, next_state => N93, 
               clocked_on => CLK_port, Q => REGISTERS_32_9_port, QN => n_2046);
   REGISTERS_reg_32_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N146, next_state => N92, 
               clocked_on => CLK_port, Q => REGISTERS_32_8_port, QN => n_2047);
   REGISTERS_reg_32_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N146, next_state => N91, 
               clocked_on => CLK_port, Q => REGISTERS_32_7_port, QN => n_2048);
   REGISTERS_reg_32_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N146, next_state => N90, 
               clocked_on => CLK_port, Q => REGISTERS_32_6_port, QN => n_2049);
   REGISTERS_reg_32_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N146, next_state => N89, 
               clocked_on => CLK_port, Q => REGISTERS_32_5_port, QN => n_2050);
   REGISTERS_reg_32_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N146, next_state => N88, 
               clocked_on => CLK_port, Q => REGISTERS_32_4_port, QN => n_2051);
   REGISTERS_reg_32_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N146, next_state => N87, 
               clocked_on => CLK_port, Q => REGISTERS_32_3_port, QN => n_2052);
   REGISTERS_reg_32_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N146, next_state => N86, 
               clocked_on => CLK_port, Q => REGISTERS_32_2_port, QN => n_2053);
   REGISTERS_reg_32_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N146, next_state => N85, 
               clocked_on => CLK_port, Q => REGISTERS_32_1_port, QN => n_2054);
   REGISTERS_reg_32_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N146, next_state => N84, 
               clocked_on => CLK_port, Q => REGISTERS_32_0_port, QN => n_2055);
   REGISTERS_reg_33_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N145, next_state => N115, 
               clocked_on => CLK_port, Q => REGISTERS_33_31_port, QN => n_2056
               );
   REGISTERS_reg_33_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N145, next_state => N114, 
               clocked_on => CLK_port, Q => REGISTERS_33_30_port, QN => n_2057
               );
   REGISTERS_reg_33_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N145, next_state => N113, 
               clocked_on => CLK_port, Q => REGISTERS_33_29_port, QN => n_2058
               );
   REGISTERS_reg_33_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N145, next_state => N112, 
               clocked_on => CLK_port, Q => REGISTERS_33_28_port, QN => n_2059
               );
   REGISTERS_reg_33_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N145, next_state => N111, 
               clocked_on => CLK_port, Q => REGISTERS_33_27_port, QN => n_2060
               );
   REGISTERS_reg_33_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N145, next_state => N110, 
               clocked_on => CLK_port, Q => REGISTERS_33_26_port, QN => n_2061
               );
   REGISTERS_reg_33_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N145, next_state => N109, 
               clocked_on => CLK_port, Q => REGISTERS_33_25_port, QN => n_2062
               );
   REGISTERS_reg_33_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N145, next_state => N108, 
               clocked_on => CLK_port, Q => REGISTERS_33_24_port, QN => n_2063
               );
   REGISTERS_reg_33_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N145, next_state => N107, 
               clocked_on => CLK_port, Q => REGISTERS_33_23_port, QN => n_2064
               );
   REGISTERS_reg_33_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N145, next_state => N106, 
               clocked_on => CLK_port, Q => REGISTERS_33_22_port, QN => n_2065
               );
   REGISTERS_reg_33_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N145, next_state => N105, 
               clocked_on => CLK_port, Q => REGISTERS_33_21_port, QN => n_2066
               );
   REGISTERS_reg_33_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N145, next_state => N104, 
               clocked_on => CLK_port, Q => REGISTERS_33_20_port, QN => n_2067
               );
   REGISTERS_reg_33_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N145, next_state => N103, 
               clocked_on => CLK_port, Q => REGISTERS_33_19_port, QN => n_2068
               );
   REGISTERS_reg_33_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N145, next_state => N102, 
               clocked_on => CLK_port, Q => REGISTERS_33_18_port, QN => n_2069
               );
   REGISTERS_reg_33_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N145, next_state => N101, 
               clocked_on => CLK_port, Q => REGISTERS_33_17_port, QN => n_2070
               );
   REGISTERS_reg_33_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N145, next_state => N100, 
               clocked_on => CLK_port, Q => REGISTERS_33_16_port, QN => n_2071
               );
   REGISTERS_reg_33_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N145, next_state => N99, 
               clocked_on => CLK_port, Q => REGISTERS_33_15_port, QN => n_2072
               );
   REGISTERS_reg_33_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N145, next_state => N98, 
               clocked_on => CLK_port, Q => REGISTERS_33_14_port, QN => n_2073
               );
   REGISTERS_reg_33_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N145, next_state => N97, 
               clocked_on => CLK_port, Q => REGISTERS_33_13_port, QN => n_2074
               );
   REGISTERS_reg_33_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N145, next_state => N96, 
               clocked_on => CLK_port, Q => REGISTERS_33_12_port, QN => n_2075
               );
   REGISTERS_reg_33_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N145, next_state => N95, 
               clocked_on => CLK_port, Q => REGISTERS_33_11_port, QN => n_2076
               );
   REGISTERS_reg_33_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N145, next_state => N94, 
               clocked_on => CLK_port, Q => REGISTERS_33_10_port, QN => n_2077
               );
   REGISTERS_reg_33_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N145, next_state => N93, 
               clocked_on => CLK_port, Q => REGISTERS_33_9_port, QN => n_2078);
   REGISTERS_reg_33_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N145, next_state => N92, 
               clocked_on => CLK_port, Q => REGISTERS_33_8_port, QN => n_2079);
   REGISTERS_reg_33_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N145, next_state => N91, 
               clocked_on => CLK_port, Q => REGISTERS_33_7_port, QN => n_2080);
   REGISTERS_reg_33_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N145, next_state => N90, 
               clocked_on => CLK_port, Q => REGISTERS_33_6_port, QN => n_2081);
   REGISTERS_reg_33_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N145, next_state => N89, 
               clocked_on => CLK_port, Q => REGISTERS_33_5_port, QN => n_2082);
   REGISTERS_reg_33_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N145, next_state => N88, 
               clocked_on => CLK_port, Q => REGISTERS_33_4_port, QN => n_2083);
   REGISTERS_reg_33_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N145, next_state => N87, 
               clocked_on => CLK_port, Q => REGISTERS_33_3_port, QN => n_2084);
   REGISTERS_reg_33_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N145, next_state => N86, 
               clocked_on => CLK_port, Q => REGISTERS_33_2_port, QN => n_2085);
   REGISTERS_reg_33_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N145, next_state => N85, 
               clocked_on => CLK_port, Q => REGISTERS_33_1_port, QN => n_2086);
   REGISTERS_reg_33_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N145, next_state => N84, 
               clocked_on => CLK_port, Q => REGISTERS_33_0_port, QN => n_2087);
   REGISTERS_reg_34_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N144, next_state => N115, 
               clocked_on => CLK_port, Q => REGISTERS_34_31_port, QN => n_2088
               );
   REGISTERS_reg_34_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N144, next_state => N114, 
               clocked_on => CLK_port, Q => REGISTERS_34_30_port, QN => n_2089
               );
   REGISTERS_reg_34_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N144, next_state => N113, 
               clocked_on => CLK_port, Q => REGISTERS_34_29_port, QN => n_2090
               );
   REGISTERS_reg_34_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N144, next_state => N112, 
               clocked_on => CLK_port, Q => REGISTERS_34_28_port, QN => n_2091
               );
   REGISTERS_reg_34_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N144, next_state => N111, 
               clocked_on => CLK_port, Q => REGISTERS_34_27_port, QN => n_2092
               );
   REGISTERS_reg_34_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N144, next_state => N110, 
               clocked_on => CLK_port, Q => REGISTERS_34_26_port, QN => n_2093
               );
   REGISTERS_reg_34_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N144, next_state => N109, 
               clocked_on => CLK_port, Q => REGISTERS_34_25_port, QN => n_2094
               );
   REGISTERS_reg_34_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N144, next_state => N108, 
               clocked_on => CLK_port, Q => REGISTERS_34_24_port, QN => n_2095
               );
   REGISTERS_reg_34_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N144, next_state => N107, 
               clocked_on => CLK_port, Q => REGISTERS_34_23_port, QN => n_2096
               );
   REGISTERS_reg_34_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N144, next_state => N106, 
               clocked_on => CLK_port, Q => REGISTERS_34_22_port, QN => n_2097
               );
   REGISTERS_reg_34_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N144, next_state => N105, 
               clocked_on => CLK_port, Q => REGISTERS_34_21_port, QN => n_2098
               );
   REGISTERS_reg_34_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N144, next_state => N104, 
               clocked_on => CLK_port, Q => REGISTERS_34_20_port, QN => n_2099
               );
   REGISTERS_reg_34_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N144, next_state => N103, 
               clocked_on => CLK_port, Q => REGISTERS_34_19_port, QN => n_2100
               );
   REGISTERS_reg_34_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N144, next_state => N102, 
               clocked_on => CLK_port, Q => REGISTERS_34_18_port, QN => n_2101
               );
   REGISTERS_reg_34_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N144, next_state => N101, 
               clocked_on => CLK_port, Q => REGISTERS_34_17_port, QN => n_2102
               );
   REGISTERS_reg_34_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N144, next_state => N100, 
               clocked_on => CLK_port, Q => REGISTERS_34_16_port, QN => n_2103
               );
   REGISTERS_reg_34_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N144, next_state => N99, 
               clocked_on => CLK_port, Q => REGISTERS_34_15_port, QN => n_2104
               );
   REGISTERS_reg_34_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N144, next_state => N98, 
               clocked_on => CLK_port, Q => REGISTERS_34_14_port, QN => n_2105
               );
   REGISTERS_reg_34_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N144, next_state => N97, 
               clocked_on => CLK_port, Q => REGISTERS_34_13_port, QN => n_2106
               );
   REGISTERS_reg_34_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N144, next_state => N96, 
               clocked_on => CLK_port, Q => REGISTERS_34_12_port, QN => n_2107
               );
   REGISTERS_reg_34_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N144, next_state => N95, 
               clocked_on => CLK_port, Q => REGISTERS_34_11_port, QN => n_2108
               );
   REGISTERS_reg_34_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N144, next_state => N94, 
               clocked_on => CLK_port, Q => REGISTERS_34_10_port, QN => n_2109
               );
   REGISTERS_reg_34_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N144, next_state => N93, 
               clocked_on => CLK_port, Q => REGISTERS_34_9_port, QN => n_2110);
   REGISTERS_reg_34_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N144, next_state => N92, 
               clocked_on => CLK_port, Q => REGISTERS_34_8_port, QN => n_2111);
   REGISTERS_reg_34_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N144, next_state => N91, 
               clocked_on => CLK_port, Q => REGISTERS_34_7_port, QN => n_2112);
   REGISTERS_reg_34_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N144, next_state => N90, 
               clocked_on => CLK_port, Q => REGISTERS_34_6_port, QN => n_2113);
   REGISTERS_reg_34_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N144, next_state => N89, 
               clocked_on => CLK_port, Q => REGISTERS_34_5_port, QN => n_2114);
   REGISTERS_reg_34_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N144, next_state => N88, 
               clocked_on => CLK_port, Q => REGISTERS_34_4_port, QN => n_2115);
   REGISTERS_reg_34_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N144, next_state => N87, 
               clocked_on => CLK_port, Q => REGISTERS_34_3_port, QN => n_2116);
   REGISTERS_reg_34_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N144, next_state => N86, 
               clocked_on => CLK_port, Q => REGISTERS_34_2_port, QN => n_2117);
   REGISTERS_reg_34_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N144, next_state => N85, 
               clocked_on => CLK_port, Q => REGISTERS_34_1_port, QN => n_2118);
   REGISTERS_reg_34_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N144, next_state => N84, 
               clocked_on => CLK_port, Q => REGISTERS_34_0_port, QN => n_2119);
   REGISTERS_reg_35_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N143, next_state => N115, 
               clocked_on => CLK_port, Q => REGISTERS_35_31_port, QN => n_2120
               );
   REGISTERS_reg_35_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N143, next_state => N114, 
               clocked_on => CLK_port, Q => REGISTERS_35_30_port, QN => n_2121
               );
   REGISTERS_reg_35_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N143, next_state => N113, 
               clocked_on => CLK_port, Q => REGISTERS_35_29_port, QN => n_2122
               );
   REGISTERS_reg_35_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N143, next_state => N112, 
               clocked_on => CLK_port, Q => REGISTERS_35_28_port, QN => n_2123
               );
   REGISTERS_reg_35_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N143, next_state => N111, 
               clocked_on => CLK_port, Q => REGISTERS_35_27_port, QN => n_2124
               );
   REGISTERS_reg_35_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N143, next_state => N110, 
               clocked_on => CLK_port, Q => REGISTERS_35_26_port, QN => n_2125
               );
   REGISTERS_reg_35_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N143, next_state => N109, 
               clocked_on => CLK_port, Q => REGISTERS_35_25_port, QN => n_2126
               );
   REGISTERS_reg_35_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N143, next_state => N108, 
               clocked_on => CLK_port, Q => REGISTERS_35_24_port, QN => n_2127
               );
   REGISTERS_reg_35_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N143, next_state => N107, 
               clocked_on => CLK_port, Q => REGISTERS_35_23_port, QN => n_2128
               );
   REGISTERS_reg_35_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N143, next_state => N106, 
               clocked_on => CLK_port, Q => REGISTERS_35_22_port, QN => n_2129
               );
   REGISTERS_reg_35_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N143, next_state => N105, 
               clocked_on => CLK_port, Q => REGISTERS_35_21_port, QN => n_2130
               );
   REGISTERS_reg_35_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N143, next_state => N104, 
               clocked_on => CLK_port, Q => REGISTERS_35_20_port, QN => n_2131
               );
   REGISTERS_reg_35_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N143, next_state => N103, 
               clocked_on => CLK_port, Q => REGISTERS_35_19_port, QN => n_2132
               );
   REGISTERS_reg_35_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N143, next_state => N102, 
               clocked_on => CLK_port, Q => REGISTERS_35_18_port, QN => n_2133
               );
   REGISTERS_reg_35_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N143, next_state => N101, 
               clocked_on => CLK_port, Q => REGISTERS_35_17_port, QN => n_2134
               );
   REGISTERS_reg_35_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N143, next_state => N100, 
               clocked_on => CLK_port, Q => REGISTERS_35_16_port, QN => n_2135
               );
   REGISTERS_reg_35_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N143, next_state => N99, 
               clocked_on => CLK_port, Q => REGISTERS_35_15_port, QN => n_2136
               );
   REGISTERS_reg_35_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N143, next_state => N98, 
               clocked_on => CLK_port, Q => REGISTERS_35_14_port, QN => n_2137
               );
   REGISTERS_reg_35_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N143, next_state => N97, 
               clocked_on => CLK_port, Q => REGISTERS_35_13_port, QN => n_2138
               );
   REGISTERS_reg_35_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N143, next_state => N96, 
               clocked_on => CLK_port, Q => REGISTERS_35_12_port, QN => n_2139
               );
   REGISTERS_reg_35_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N143, next_state => N95, 
               clocked_on => CLK_port, Q => REGISTERS_35_11_port, QN => n_2140
               );
   REGISTERS_reg_35_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N143, next_state => N94, 
               clocked_on => CLK_port, Q => REGISTERS_35_10_port, QN => n_2141
               );
   REGISTERS_reg_35_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N143, next_state => N93, 
               clocked_on => CLK_port, Q => REGISTERS_35_9_port, QN => n_2142);
   REGISTERS_reg_35_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N143, next_state => N92, 
               clocked_on => CLK_port, Q => REGISTERS_35_8_port, QN => n_2143);
   REGISTERS_reg_35_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N143, next_state => N91, 
               clocked_on => CLK_port, Q => REGISTERS_35_7_port, QN => n_2144);
   REGISTERS_reg_35_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N143, next_state => N90, 
               clocked_on => CLK_port, Q => REGISTERS_35_6_port, QN => n_2145);
   REGISTERS_reg_35_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N143, next_state => N89, 
               clocked_on => CLK_port, Q => REGISTERS_35_5_port, QN => n_2146);
   REGISTERS_reg_35_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N143, next_state => N88, 
               clocked_on => CLK_port, Q => REGISTERS_35_4_port, QN => n_2147);
   REGISTERS_reg_35_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N143, next_state => N87, 
               clocked_on => CLK_port, Q => REGISTERS_35_3_port, QN => n_2148);
   REGISTERS_reg_35_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N143, next_state => N86, 
               clocked_on => CLK_port, Q => REGISTERS_35_2_port, QN => n_2149);
   REGISTERS_reg_35_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N143, next_state => N85, 
               clocked_on => CLK_port, Q => REGISTERS_35_1_port, QN => n_2150);
   REGISTERS_reg_35_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N143, next_state => N84, 
               clocked_on => CLK_port, Q => REGISTERS_35_0_port, QN => n_2151);
   REGISTERS_reg_36_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N142, next_state => N115, 
               clocked_on => CLK_port, Q => REGISTERS_36_31_port, QN => n_2152
               );
   REGISTERS_reg_36_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N142, next_state => N114, 
               clocked_on => CLK_port, Q => REGISTERS_36_30_port, QN => n_2153
               );
   REGISTERS_reg_36_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N142, next_state => N113, 
               clocked_on => CLK_port, Q => REGISTERS_36_29_port, QN => n_2154
               );
   REGISTERS_reg_36_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N142, next_state => N112, 
               clocked_on => CLK_port, Q => REGISTERS_36_28_port, QN => n_2155
               );
   REGISTERS_reg_36_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N142, next_state => N111, 
               clocked_on => CLK_port, Q => REGISTERS_36_27_port, QN => n_2156
               );
   REGISTERS_reg_36_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N142, next_state => N110, 
               clocked_on => CLK_port, Q => REGISTERS_36_26_port, QN => n_2157
               );
   REGISTERS_reg_36_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N142, next_state => N109, 
               clocked_on => CLK_port, Q => REGISTERS_36_25_port, QN => n_2158
               );
   REGISTERS_reg_36_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N142, next_state => N108, 
               clocked_on => CLK_port, Q => REGISTERS_36_24_port, QN => n_2159
               );
   REGISTERS_reg_36_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N142, next_state => N107, 
               clocked_on => CLK_port, Q => REGISTERS_36_23_port, QN => n_2160
               );
   REGISTERS_reg_36_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N142, next_state => N106, 
               clocked_on => CLK_port, Q => REGISTERS_36_22_port, QN => n_2161
               );
   REGISTERS_reg_36_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N142, next_state => N105, 
               clocked_on => CLK_port, Q => REGISTERS_36_21_port, QN => n_2162
               );
   REGISTERS_reg_36_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N142, next_state => N104, 
               clocked_on => CLK_port, Q => REGISTERS_36_20_port, QN => n_2163
               );
   REGISTERS_reg_36_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N142, next_state => N103, 
               clocked_on => CLK_port, Q => REGISTERS_36_19_port, QN => n_2164
               );
   REGISTERS_reg_36_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N142, next_state => N102, 
               clocked_on => CLK_port, Q => REGISTERS_36_18_port, QN => n_2165
               );
   REGISTERS_reg_36_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N142, next_state => N101, 
               clocked_on => CLK_port, Q => REGISTERS_36_17_port, QN => n_2166
               );
   REGISTERS_reg_36_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N142, next_state => N100, 
               clocked_on => CLK_port, Q => REGISTERS_36_16_port, QN => n_2167
               );
   REGISTERS_reg_36_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N142, next_state => N99, 
               clocked_on => CLK_port, Q => REGISTERS_36_15_port, QN => n_2168
               );
   REGISTERS_reg_36_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N142, next_state => N98, 
               clocked_on => CLK_port, Q => REGISTERS_36_14_port, QN => n_2169
               );
   REGISTERS_reg_36_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N142, next_state => N97, 
               clocked_on => CLK_port, Q => REGISTERS_36_13_port, QN => n_2170
               );
   REGISTERS_reg_36_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N142, next_state => N96, 
               clocked_on => CLK_port, Q => REGISTERS_36_12_port, QN => n_2171
               );
   REGISTERS_reg_36_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N142, next_state => N95, 
               clocked_on => CLK_port, Q => REGISTERS_36_11_port, QN => n_2172
               );
   REGISTERS_reg_36_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N142, next_state => N94, 
               clocked_on => CLK_port, Q => REGISTERS_36_10_port, QN => n_2173
               );
   REGISTERS_reg_36_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N142, next_state => N93, 
               clocked_on => CLK_port, Q => REGISTERS_36_9_port, QN => n_2174);
   REGISTERS_reg_36_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N142, next_state => N92, 
               clocked_on => CLK_port, Q => REGISTERS_36_8_port, QN => n_2175);
   REGISTERS_reg_36_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N142, next_state => N91, 
               clocked_on => CLK_port, Q => REGISTERS_36_7_port, QN => n_2176);
   REGISTERS_reg_36_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N142, next_state => N90, 
               clocked_on => CLK_port, Q => REGISTERS_36_6_port, QN => n_2177);
   REGISTERS_reg_36_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N142, next_state => N89, 
               clocked_on => CLK_port, Q => REGISTERS_36_5_port, QN => n_2178);
   REGISTERS_reg_36_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N142, next_state => N88, 
               clocked_on => CLK_port, Q => REGISTERS_36_4_port, QN => n_2179);
   REGISTERS_reg_36_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N142, next_state => N87, 
               clocked_on => CLK_port, Q => REGISTERS_36_3_port, QN => n_2180);
   REGISTERS_reg_36_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N142, next_state => N86, 
               clocked_on => CLK_port, Q => REGISTERS_36_2_port, QN => n_2181);
   REGISTERS_reg_36_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N142, next_state => N85, 
               clocked_on => CLK_port, Q => REGISTERS_36_1_port, QN => n_2182);
   REGISTERS_reg_36_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N142, next_state => N84, 
               clocked_on => CLK_port, Q => REGISTERS_36_0_port, QN => n_2183);
   REGISTERS_reg_37_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N141, next_state => N115, 
               clocked_on => CLK_port, Q => REGISTERS_37_31_port, QN => n_2184
               );
   REGISTERS_reg_37_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N141, next_state => N114, 
               clocked_on => CLK_port, Q => REGISTERS_37_30_port, QN => n_2185
               );
   REGISTERS_reg_37_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N141, next_state => N113, 
               clocked_on => CLK_port, Q => REGISTERS_37_29_port, QN => n_2186
               );
   REGISTERS_reg_37_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N141, next_state => N112, 
               clocked_on => CLK_port, Q => REGISTERS_37_28_port, QN => n_2187
               );
   REGISTERS_reg_37_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N141, next_state => N111, 
               clocked_on => CLK_port, Q => REGISTERS_37_27_port, QN => n_2188
               );
   REGISTERS_reg_37_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N141, next_state => N110, 
               clocked_on => CLK_port, Q => REGISTERS_37_26_port, QN => n_2189
               );
   REGISTERS_reg_37_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N141, next_state => N109, 
               clocked_on => CLK_port, Q => REGISTERS_37_25_port, QN => n_2190
               );
   REGISTERS_reg_37_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N141, next_state => N108, 
               clocked_on => CLK_port, Q => REGISTERS_37_24_port, QN => n_2191
               );
   REGISTERS_reg_37_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N141, next_state => N107, 
               clocked_on => CLK_port, Q => REGISTERS_37_23_port, QN => n_2192
               );
   REGISTERS_reg_37_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N141, next_state => N106, 
               clocked_on => CLK_port, Q => REGISTERS_37_22_port, QN => n_2193
               );
   REGISTERS_reg_37_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N141, next_state => N105, 
               clocked_on => CLK_port, Q => REGISTERS_37_21_port, QN => n_2194
               );
   REGISTERS_reg_37_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N141, next_state => N104, 
               clocked_on => CLK_port, Q => REGISTERS_37_20_port, QN => n_2195
               );
   REGISTERS_reg_37_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N141, next_state => N103, 
               clocked_on => CLK_port, Q => REGISTERS_37_19_port, QN => n_2196
               );
   REGISTERS_reg_37_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N141, next_state => N102, 
               clocked_on => CLK_port, Q => REGISTERS_37_18_port, QN => n_2197
               );
   REGISTERS_reg_37_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N141, next_state => N101, 
               clocked_on => CLK_port, Q => REGISTERS_37_17_port, QN => n_2198
               );
   REGISTERS_reg_37_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N141, next_state => N100, 
               clocked_on => CLK_port, Q => REGISTERS_37_16_port, QN => n_2199
               );
   REGISTERS_reg_37_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N141, next_state => N99, 
               clocked_on => CLK_port, Q => REGISTERS_37_15_port, QN => n_2200
               );
   REGISTERS_reg_37_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N141, next_state => N98, 
               clocked_on => CLK_port, Q => REGISTERS_37_14_port, QN => n_2201
               );
   REGISTERS_reg_37_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N141, next_state => N97, 
               clocked_on => CLK_port, Q => REGISTERS_37_13_port, QN => n_2202
               );
   REGISTERS_reg_37_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N141, next_state => N96, 
               clocked_on => CLK_port, Q => REGISTERS_37_12_port, QN => n_2203
               );
   REGISTERS_reg_37_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N141, next_state => N95, 
               clocked_on => CLK_port, Q => REGISTERS_37_11_port, QN => n_2204
               );
   REGISTERS_reg_37_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N141, next_state => N94, 
               clocked_on => CLK_port, Q => REGISTERS_37_10_port, QN => n_2205
               );
   REGISTERS_reg_37_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N141, next_state => N93, 
               clocked_on => CLK_port, Q => REGISTERS_37_9_port, QN => n_2206);
   REGISTERS_reg_37_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N141, next_state => N92, 
               clocked_on => CLK_port, Q => REGISTERS_37_8_port, QN => n_2207);
   REGISTERS_reg_37_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N141, next_state => N91, 
               clocked_on => CLK_port, Q => REGISTERS_37_7_port, QN => n_2208);
   REGISTERS_reg_37_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N141, next_state => N90, 
               clocked_on => CLK_port, Q => REGISTERS_37_6_port, QN => n_2209);
   REGISTERS_reg_37_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N141, next_state => N89, 
               clocked_on => CLK_port, Q => REGISTERS_37_5_port, QN => n_2210);
   REGISTERS_reg_37_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N141, next_state => N88, 
               clocked_on => CLK_port, Q => REGISTERS_37_4_port, QN => n_2211);
   REGISTERS_reg_37_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N141, next_state => N87, 
               clocked_on => CLK_port, Q => REGISTERS_37_3_port, QN => n_2212);
   REGISTERS_reg_37_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N141, next_state => N86, 
               clocked_on => CLK_port, Q => REGISTERS_37_2_port, QN => n_2213);
   REGISTERS_reg_37_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N141, next_state => N85, 
               clocked_on => CLK_port, Q => REGISTERS_37_1_port, QN => n_2214);
   REGISTERS_reg_37_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N141, next_state => N84, 
               clocked_on => CLK_port, Q => REGISTERS_37_0_port, QN => n_2215);
   REGISTERS_reg_38_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N140, next_state => N115, 
               clocked_on => CLK_port, Q => REGISTERS_38_31_port, QN => n_2216
               );
   REGISTERS_reg_38_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N140, next_state => N114, 
               clocked_on => CLK_port, Q => REGISTERS_38_30_port, QN => n_2217
               );
   REGISTERS_reg_38_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N140, next_state => N113, 
               clocked_on => CLK_port, Q => REGISTERS_38_29_port, QN => n_2218
               );
   REGISTERS_reg_38_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N140, next_state => N112, 
               clocked_on => CLK_port, Q => REGISTERS_38_28_port, QN => n_2219
               );
   REGISTERS_reg_38_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N140, next_state => N111, 
               clocked_on => CLK_port, Q => REGISTERS_38_27_port, QN => n_2220
               );
   REGISTERS_reg_38_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N140, next_state => N110, 
               clocked_on => CLK_port, Q => REGISTERS_38_26_port, QN => n_2221
               );
   REGISTERS_reg_38_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N140, next_state => N109, 
               clocked_on => CLK_port, Q => REGISTERS_38_25_port, QN => n_2222
               );
   REGISTERS_reg_38_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N140, next_state => N108, 
               clocked_on => CLK_port, Q => REGISTERS_38_24_port, QN => n_2223
               );
   REGISTERS_reg_38_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N140, next_state => N107, 
               clocked_on => CLK_port, Q => REGISTERS_38_23_port, QN => n_2224
               );
   REGISTERS_reg_38_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N140, next_state => N106, 
               clocked_on => CLK_port, Q => REGISTERS_38_22_port, QN => n_2225
               );
   REGISTERS_reg_38_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N140, next_state => N105, 
               clocked_on => CLK_port, Q => REGISTERS_38_21_port, QN => n_2226
               );
   REGISTERS_reg_38_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N140, next_state => N104, 
               clocked_on => CLK_port, Q => REGISTERS_38_20_port, QN => n_2227
               );
   REGISTERS_reg_38_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N140, next_state => N103, 
               clocked_on => CLK_port, Q => REGISTERS_38_19_port, QN => n_2228
               );
   REGISTERS_reg_38_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N140, next_state => N102, 
               clocked_on => CLK_port, Q => REGISTERS_38_18_port, QN => n_2229
               );
   REGISTERS_reg_38_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N140, next_state => N101, 
               clocked_on => CLK_port, Q => REGISTERS_38_17_port, QN => n_2230
               );
   REGISTERS_reg_38_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N140, next_state => N100, 
               clocked_on => CLK_port, Q => REGISTERS_38_16_port, QN => n_2231
               );
   REGISTERS_reg_38_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N140, next_state => N99, 
               clocked_on => CLK_port, Q => REGISTERS_38_15_port, QN => n_2232
               );
   REGISTERS_reg_38_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N140, next_state => N98, 
               clocked_on => CLK_port, Q => REGISTERS_38_14_port, QN => n_2233
               );
   REGISTERS_reg_38_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N140, next_state => N97, 
               clocked_on => CLK_port, Q => REGISTERS_38_13_port, QN => n_2234
               );
   REGISTERS_reg_38_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N140, next_state => N96, 
               clocked_on => CLK_port, Q => REGISTERS_38_12_port, QN => n_2235
               );
   REGISTERS_reg_38_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N140, next_state => N95, 
               clocked_on => CLK_port, Q => REGISTERS_38_11_port, QN => n_2236
               );
   REGISTERS_reg_38_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N140, next_state => N94, 
               clocked_on => CLK_port, Q => REGISTERS_38_10_port, QN => n_2237
               );
   REGISTERS_reg_38_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N140, next_state => N93, 
               clocked_on => CLK_port, Q => REGISTERS_38_9_port, QN => n_2238);
   REGISTERS_reg_38_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N140, next_state => N92, 
               clocked_on => CLK_port, Q => REGISTERS_38_8_port, QN => n_2239);
   REGISTERS_reg_38_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N140, next_state => N91, 
               clocked_on => CLK_port, Q => REGISTERS_38_7_port, QN => n_2240);
   REGISTERS_reg_38_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N140, next_state => N90, 
               clocked_on => CLK_port, Q => REGISTERS_38_6_port, QN => n_2241);
   REGISTERS_reg_38_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N140, next_state => N89, 
               clocked_on => CLK_port, Q => REGISTERS_38_5_port, QN => n_2242);
   REGISTERS_reg_38_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N140, next_state => N88, 
               clocked_on => CLK_port, Q => REGISTERS_38_4_port, QN => n_2243);
   REGISTERS_reg_38_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N140, next_state => N87, 
               clocked_on => CLK_port, Q => REGISTERS_38_3_port, QN => n_2244);
   REGISTERS_reg_38_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N140, next_state => N86, 
               clocked_on => CLK_port, Q => REGISTERS_38_2_port, QN => n_2245);
   REGISTERS_reg_38_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N140, next_state => N85, 
               clocked_on => CLK_port, Q => REGISTERS_38_1_port, QN => n_2246);
   REGISTERS_reg_38_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N140, next_state => N84, 
               clocked_on => CLK_port, Q => REGISTERS_38_0_port, QN => n_2247);
   REGISTERS_reg_39_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N139, next_state => N115, 
               clocked_on => CLK_port, Q => REGISTERS_39_31_port, QN => n_2248
               );
   REGISTERS_reg_39_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N139, next_state => N114, 
               clocked_on => CLK_port, Q => REGISTERS_39_30_port, QN => n_2249
               );
   REGISTERS_reg_39_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N139, next_state => N113, 
               clocked_on => CLK_port, Q => REGISTERS_39_29_port, QN => n_2250
               );
   REGISTERS_reg_39_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N139, next_state => N112, 
               clocked_on => CLK_port, Q => REGISTERS_39_28_port, QN => n_2251
               );
   REGISTERS_reg_39_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N139, next_state => N111, 
               clocked_on => CLK_port, Q => REGISTERS_39_27_port, QN => n_2252
               );
   REGISTERS_reg_39_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N139, next_state => N110, 
               clocked_on => CLK_port, Q => REGISTERS_39_26_port, QN => n_2253
               );
   REGISTERS_reg_39_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N139, next_state => N109, 
               clocked_on => CLK_port, Q => REGISTERS_39_25_port, QN => n_2254
               );
   REGISTERS_reg_39_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N139, next_state => N108, 
               clocked_on => CLK_port, Q => REGISTERS_39_24_port, QN => n_2255
               );
   REGISTERS_reg_39_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N139, next_state => N107, 
               clocked_on => CLK_port, Q => REGISTERS_39_23_port, QN => n_2256
               );
   REGISTERS_reg_39_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N139, next_state => N106, 
               clocked_on => CLK_port, Q => REGISTERS_39_22_port, QN => n_2257
               );
   REGISTERS_reg_39_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N139, next_state => N105, 
               clocked_on => CLK_port, Q => REGISTERS_39_21_port, QN => n_2258
               );
   REGISTERS_reg_39_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N139, next_state => N104, 
               clocked_on => CLK_port, Q => REGISTERS_39_20_port, QN => n_2259
               );
   REGISTERS_reg_39_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N139, next_state => N103, 
               clocked_on => CLK_port, Q => REGISTERS_39_19_port, QN => n_2260
               );
   REGISTERS_reg_39_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N139, next_state => N102, 
               clocked_on => CLK_port, Q => REGISTERS_39_18_port, QN => n_2261
               );
   REGISTERS_reg_39_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N139, next_state => N101, 
               clocked_on => CLK_port, Q => REGISTERS_39_17_port, QN => n_2262
               );
   REGISTERS_reg_39_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N139, next_state => N100, 
               clocked_on => CLK_port, Q => REGISTERS_39_16_port, QN => n_2263
               );
   REGISTERS_reg_39_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N139, next_state => N99, 
               clocked_on => CLK_port, Q => REGISTERS_39_15_port, QN => n_2264
               );
   REGISTERS_reg_39_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N139, next_state => N98, 
               clocked_on => CLK_port, Q => REGISTERS_39_14_port, QN => n_2265
               );
   REGISTERS_reg_39_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N139, next_state => N97, 
               clocked_on => CLK_port, Q => REGISTERS_39_13_port, QN => n_2266
               );
   REGISTERS_reg_39_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N139, next_state => N96, 
               clocked_on => CLK_port, Q => REGISTERS_39_12_port, QN => n_2267
               );
   REGISTERS_reg_39_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N139, next_state => N95, 
               clocked_on => CLK_port, Q => REGISTERS_39_11_port, QN => n_2268
               );
   REGISTERS_reg_39_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N139, next_state => N94, 
               clocked_on => CLK_port, Q => REGISTERS_39_10_port, QN => n_2269
               );
   REGISTERS_reg_39_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N139, next_state => N93, 
               clocked_on => CLK_port, Q => REGISTERS_39_9_port, QN => n_2270);
   REGISTERS_reg_39_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N139, next_state => N92, 
               clocked_on => CLK_port, Q => REGISTERS_39_8_port, QN => n_2271);
   REGISTERS_reg_39_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N139, next_state => N91, 
               clocked_on => CLK_port, Q => REGISTERS_39_7_port, QN => n_2272);
   REGISTERS_reg_39_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N139, next_state => N90, 
               clocked_on => CLK_port, Q => REGISTERS_39_6_port, QN => n_2273);
   REGISTERS_reg_39_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N139, next_state => N89, 
               clocked_on => CLK_port, Q => REGISTERS_39_5_port, QN => n_2274);
   REGISTERS_reg_39_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N139, next_state => N88, 
               clocked_on => CLK_port, Q => REGISTERS_39_4_port, QN => n_2275);
   REGISTERS_reg_39_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N139, next_state => N87, 
               clocked_on => CLK_port, Q => REGISTERS_39_3_port, QN => n_2276);
   REGISTERS_reg_39_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N139, next_state => N86, 
               clocked_on => CLK_port, Q => REGISTERS_39_2_port, QN => n_2277);
   REGISTERS_reg_39_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N139, next_state => N85, 
               clocked_on => CLK_port, Q => REGISTERS_39_1_port, QN => n_2278);
   REGISTERS_reg_39_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N139, next_state => N84, 
               clocked_on => CLK_port, Q => REGISTERS_39_0_port, QN => n_2279);
   REGISTERS_reg_40_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N138, next_state => N115, 
               clocked_on => CLK_port, Q => REGISTERS_40_31_port, QN => n_2280
               );
   REGISTERS_reg_40_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N138, next_state => N114, 
               clocked_on => CLK_port, Q => REGISTERS_40_30_port, QN => n_2281
               );
   REGISTERS_reg_40_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N138, next_state => N113, 
               clocked_on => CLK_port, Q => REGISTERS_40_29_port, QN => n_2282
               );
   REGISTERS_reg_40_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N138, next_state => N112, 
               clocked_on => CLK_port, Q => REGISTERS_40_28_port, QN => n_2283
               );
   REGISTERS_reg_40_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N138, next_state => N111, 
               clocked_on => CLK_port, Q => REGISTERS_40_27_port, QN => n_2284
               );
   REGISTERS_reg_40_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N138, next_state => N110, 
               clocked_on => CLK_port, Q => REGISTERS_40_26_port, QN => n_2285
               );
   REGISTERS_reg_40_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N138, next_state => N109, 
               clocked_on => CLK_port, Q => REGISTERS_40_25_port, QN => n_2286
               );
   REGISTERS_reg_40_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N138, next_state => N108, 
               clocked_on => CLK_port, Q => REGISTERS_40_24_port, QN => n_2287
               );
   REGISTERS_reg_40_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N138, next_state => N107, 
               clocked_on => CLK_port, Q => REGISTERS_40_23_port, QN => n_2288
               );
   REGISTERS_reg_40_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N138, next_state => N106, 
               clocked_on => CLK_port, Q => REGISTERS_40_22_port, QN => n_2289
               );
   REGISTERS_reg_40_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N138, next_state => N105, 
               clocked_on => CLK_port, Q => REGISTERS_40_21_port, QN => n_2290
               );
   REGISTERS_reg_40_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N138, next_state => N104, 
               clocked_on => CLK_port, Q => REGISTERS_40_20_port, QN => n_2291
               );
   REGISTERS_reg_40_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N138, next_state => N103, 
               clocked_on => CLK_port, Q => REGISTERS_40_19_port, QN => n_2292
               );
   REGISTERS_reg_40_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N138, next_state => N102, 
               clocked_on => CLK_port, Q => REGISTERS_40_18_port, QN => n_2293
               );
   REGISTERS_reg_40_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N138, next_state => N101, 
               clocked_on => CLK_port, Q => REGISTERS_40_17_port, QN => n_2294
               );
   REGISTERS_reg_40_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N138, next_state => N100, 
               clocked_on => CLK_port, Q => REGISTERS_40_16_port, QN => n_2295
               );
   REGISTERS_reg_40_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N138, next_state => N99, 
               clocked_on => CLK_port, Q => REGISTERS_40_15_port, QN => n_2296
               );
   REGISTERS_reg_40_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N138, next_state => N98, 
               clocked_on => CLK_port, Q => REGISTERS_40_14_port, QN => n_2297
               );
   REGISTERS_reg_40_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N138, next_state => N97, 
               clocked_on => CLK_port, Q => REGISTERS_40_13_port, QN => n_2298
               );
   REGISTERS_reg_40_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N138, next_state => N96, 
               clocked_on => CLK_port, Q => REGISTERS_40_12_port, QN => n_2299
               );
   REGISTERS_reg_40_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N138, next_state => N95, 
               clocked_on => CLK_port, Q => REGISTERS_40_11_port, QN => n_2300
               );
   REGISTERS_reg_40_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N138, next_state => N94, 
               clocked_on => CLK_port, Q => REGISTERS_40_10_port, QN => n_2301
               );
   REGISTERS_reg_40_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N138, next_state => N93, 
               clocked_on => CLK_port, Q => REGISTERS_40_9_port, QN => n_2302);
   REGISTERS_reg_40_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N138, next_state => N92, 
               clocked_on => CLK_port, Q => REGISTERS_40_8_port, QN => n_2303);
   REGISTERS_reg_40_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N138, next_state => N91, 
               clocked_on => CLK_port, Q => REGISTERS_40_7_port, QN => n_2304);
   REGISTERS_reg_40_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N138, next_state => N90, 
               clocked_on => CLK_port, Q => REGISTERS_40_6_port, QN => n_2305);
   REGISTERS_reg_40_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N138, next_state => N89, 
               clocked_on => CLK_port, Q => REGISTERS_40_5_port, QN => n_2306);
   REGISTERS_reg_40_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N138, next_state => N88, 
               clocked_on => CLK_port, Q => REGISTERS_40_4_port, QN => n_2307);
   REGISTERS_reg_40_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N138, next_state => N87, 
               clocked_on => CLK_port, Q => REGISTERS_40_3_port, QN => n_2308);
   REGISTERS_reg_40_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N138, next_state => N86, 
               clocked_on => CLK_port, Q => REGISTERS_40_2_port, QN => n_2309);
   REGISTERS_reg_40_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N138, next_state => N85, 
               clocked_on => CLK_port, Q => REGISTERS_40_1_port, QN => n_2310);
   REGISTERS_reg_40_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N138, next_state => N84, 
               clocked_on => CLK_port, Q => REGISTERS_40_0_port, QN => n_2311);
   REGISTERS_reg_41_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N137, next_state => N115, 
               clocked_on => CLK_port, Q => REGISTERS_41_31_port, QN => n_2312
               );
   REGISTERS_reg_41_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N137, next_state => N114, 
               clocked_on => CLK_port, Q => REGISTERS_41_30_port, QN => n_2313
               );
   REGISTERS_reg_41_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N137, next_state => N113, 
               clocked_on => CLK_port, Q => REGISTERS_41_29_port, QN => n_2314
               );
   REGISTERS_reg_41_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N137, next_state => N112, 
               clocked_on => CLK_port, Q => REGISTERS_41_28_port, QN => n_2315
               );
   REGISTERS_reg_41_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N137, next_state => N111, 
               clocked_on => CLK_port, Q => REGISTERS_41_27_port, QN => n_2316
               );
   REGISTERS_reg_41_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N137, next_state => N110, 
               clocked_on => CLK_port, Q => REGISTERS_41_26_port, QN => n_2317
               );
   REGISTERS_reg_41_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N137, next_state => N109, 
               clocked_on => CLK_port, Q => REGISTERS_41_25_port, QN => n_2318
               );
   REGISTERS_reg_41_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N137, next_state => N108, 
               clocked_on => CLK_port, Q => REGISTERS_41_24_port, QN => n_2319
               );
   REGISTERS_reg_41_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N137, next_state => N107, 
               clocked_on => CLK_port, Q => REGISTERS_41_23_port, QN => n_2320
               );
   REGISTERS_reg_41_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N137, next_state => N106, 
               clocked_on => CLK_port, Q => REGISTERS_41_22_port, QN => n_2321
               );
   REGISTERS_reg_41_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N137, next_state => N105, 
               clocked_on => CLK_port, Q => REGISTERS_41_21_port, QN => n_2322
               );
   REGISTERS_reg_41_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N137, next_state => N104, 
               clocked_on => CLK_port, Q => REGISTERS_41_20_port, QN => n_2323
               );
   REGISTERS_reg_41_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N137, next_state => N103, 
               clocked_on => CLK_port, Q => REGISTERS_41_19_port, QN => n_2324
               );
   REGISTERS_reg_41_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N137, next_state => N102, 
               clocked_on => CLK_port, Q => REGISTERS_41_18_port, QN => n_2325
               );
   REGISTERS_reg_41_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N137, next_state => N101, 
               clocked_on => CLK_port, Q => REGISTERS_41_17_port, QN => n_2326
               );
   REGISTERS_reg_41_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N137, next_state => N100, 
               clocked_on => CLK_port, Q => REGISTERS_41_16_port, QN => n_2327
               );
   REGISTERS_reg_41_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N137, next_state => N99, 
               clocked_on => CLK_port, Q => REGISTERS_41_15_port, QN => n_2328
               );
   REGISTERS_reg_41_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N137, next_state => N98, 
               clocked_on => CLK_port, Q => REGISTERS_41_14_port, QN => n_2329
               );
   REGISTERS_reg_41_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N137, next_state => N97, 
               clocked_on => CLK_port, Q => REGISTERS_41_13_port, QN => n_2330
               );
   REGISTERS_reg_41_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N137, next_state => N96, 
               clocked_on => CLK_port, Q => REGISTERS_41_12_port, QN => n_2331
               );
   REGISTERS_reg_41_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N137, next_state => N95, 
               clocked_on => CLK_port, Q => REGISTERS_41_11_port, QN => n_2332
               );
   REGISTERS_reg_41_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N137, next_state => N94, 
               clocked_on => CLK_port, Q => REGISTERS_41_10_port, QN => n_2333
               );
   REGISTERS_reg_41_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N137, next_state => N93, 
               clocked_on => CLK_port, Q => REGISTERS_41_9_port, QN => n_2334);
   REGISTERS_reg_41_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N137, next_state => N92, 
               clocked_on => CLK_port, Q => REGISTERS_41_8_port, QN => n_2335);
   REGISTERS_reg_41_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N137, next_state => N91, 
               clocked_on => CLK_port, Q => REGISTERS_41_7_port, QN => n_2336);
   REGISTERS_reg_41_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N137, next_state => N90, 
               clocked_on => CLK_port, Q => REGISTERS_41_6_port, QN => n_2337);
   REGISTERS_reg_41_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N137, next_state => N89, 
               clocked_on => CLK_port, Q => REGISTERS_41_5_port, QN => n_2338);
   REGISTERS_reg_41_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N137, next_state => N88, 
               clocked_on => CLK_port, Q => REGISTERS_41_4_port, QN => n_2339);
   REGISTERS_reg_41_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N137, next_state => N87, 
               clocked_on => CLK_port, Q => REGISTERS_41_3_port, QN => n_2340);
   REGISTERS_reg_41_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N137, next_state => N86, 
               clocked_on => CLK_port, Q => REGISTERS_41_2_port, QN => n_2341);
   REGISTERS_reg_41_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N137, next_state => N85, 
               clocked_on => CLK_port, Q => REGISTERS_41_1_port, QN => n_2342);
   REGISTERS_reg_41_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N137, next_state => N84, 
               clocked_on => CLK_port, Q => REGISTERS_41_0_port, QN => n_2343);
   REGISTERS_reg_42_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N136, next_state => N115, 
               clocked_on => CLK_port, Q => REGISTERS_42_31_port, QN => n_2344
               );
   REGISTERS_reg_42_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N136, next_state => N114, 
               clocked_on => CLK_port, Q => REGISTERS_42_30_port, QN => n_2345
               );
   REGISTERS_reg_42_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N136, next_state => N113, 
               clocked_on => CLK_port, Q => REGISTERS_42_29_port, QN => n_2346
               );
   REGISTERS_reg_42_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N136, next_state => N112, 
               clocked_on => CLK_port, Q => REGISTERS_42_28_port, QN => n_2347
               );
   REGISTERS_reg_42_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N136, next_state => N111, 
               clocked_on => CLK_port, Q => REGISTERS_42_27_port, QN => n_2348
               );
   REGISTERS_reg_42_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N136, next_state => N110, 
               clocked_on => CLK_port, Q => REGISTERS_42_26_port, QN => n_2349
               );
   REGISTERS_reg_42_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N136, next_state => N109, 
               clocked_on => CLK_port, Q => REGISTERS_42_25_port, QN => n_2350
               );
   REGISTERS_reg_42_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N136, next_state => N108, 
               clocked_on => CLK_port, Q => REGISTERS_42_24_port, QN => n_2351
               );
   REGISTERS_reg_42_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N136, next_state => N107, 
               clocked_on => CLK_port, Q => REGISTERS_42_23_port, QN => n_2352
               );
   REGISTERS_reg_42_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N136, next_state => N106, 
               clocked_on => CLK_port, Q => REGISTERS_42_22_port, QN => n_2353
               );
   REGISTERS_reg_42_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N136, next_state => N105, 
               clocked_on => CLK_port, Q => REGISTERS_42_21_port, QN => n_2354
               );
   REGISTERS_reg_42_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N136, next_state => N104, 
               clocked_on => CLK_port, Q => REGISTERS_42_20_port, QN => n_2355
               );
   REGISTERS_reg_42_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N136, next_state => N103, 
               clocked_on => CLK_port, Q => REGISTERS_42_19_port, QN => n_2356
               );
   REGISTERS_reg_42_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N136, next_state => N102, 
               clocked_on => CLK_port, Q => REGISTERS_42_18_port, QN => n_2357
               );
   REGISTERS_reg_42_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N136, next_state => N101, 
               clocked_on => CLK_port, Q => REGISTERS_42_17_port, QN => n_2358
               );
   REGISTERS_reg_42_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N136, next_state => N100, 
               clocked_on => CLK_port, Q => REGISTERS_42_16_port, QN => n_2359
               );
   REGISTERS_reg_42_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N136, next_state => N99, 
               clocked_on => CLK_port, Q => REGISTERS_42_15_port, QN => n_2360
               );
   REGISTERS_reg_42_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N136, next_state => N98, 
               clocked_on => CLK_port, Q => REGISTERS_42_14_port, QN => n_2361
               );
   REGISTERS_reg_42_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N136, next_state => N97, 
               clocked_on => CLK_port, Q => REGISTERS_42_13_port, QN => n_2362
               );
   REGISTERS_reg_42_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N136, next_state => N96, 
               clocked_on => CLK_port, Q => REGISTERS_42_12_port, QN => n_2363
               );
   REGISTERS_reg_42_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N136, next_state => N95, 
               clocked_on => CLK_port, Q => REGISTERS_42_11_port, QN => n_2364
               );
   REGISTERS_reg_42_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N136, next_state => N94, 
               clocked_on => CLK_port, Q => REGISTERS_42_10_port, QN => n_2365
               );
   REGISTERS_reg_42_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N136, next_state => N93, 
               clocked_on => CLK_port, Q => REGISTERS_42_9_port, QN => n_2366);
   REGISTERS_reg_42_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N136, next_state => N92, 
               clocked_on => CLK_port, Q => REGISTERS_42_8_port, QN => n_2367);
   REGISTERS_reg_42_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N136, next_state => N91, 
               clocked_on => CLK_port, Q => REGISTERS_42_7_port, QN => n_2368);
   REGISTERS_reg_42_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N136, next_state => N90, 
               clocked_on => CLK_port, Q => REGISTERS_42_6_port, QN => n_2369);
   REGISTERS_reg_42_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N136, next_state => N89, 
               clocked_on => CLK_port, Q => REGISTERS_42_5_port, QN => n_2370);
   REGISTERS_reg_42_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N136, next_state => N88, 
               clocked_on => CLK_port, Q => REGISTERS_42_4_port, QN => n_2371);
   REGISTERS_reg_42_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N136, next_state => N87, 
               clocked_on => CLK_port, Q => REGISTERS_42_3_port, QN => n_2372);
   REGISTERS_reg_42_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N136, next_state => N86, 
               clocked_on => CLK_port, Q => REGISTERS_42_2_port, QN => n_2373);
   REGISTERS_reg_42_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N136, next_state => N85, 
               clocked_on => CLK_port, Q => REGISTERS_42_1_port, QN => n_2374);
   REGISTERS_reg_42_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N136, next_state => N84, 
               clocked_on => CLK_port, Q => REGISTERS_42_0_port, QN => n_2375);
   REGISTERS_reg_43_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N135, next_state => N115, 
               clocked_on => CLK_port, Q => REGISTERS_43_31_port, QN => n_2376
               );
   REGISTERS_reg_43_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N135, next_state => N114, 
               clocked_on => CLK_port, Q => REGISTERS_43_30_port, QN => n_2377
               );
   REGISTERS_reg_43_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N135, next_state => N113, 
               clocked_on => CLK_port, Q => REGISTERS_43_29_port, QN => n_2378
               );
   REGISTERS_reg_43_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N135, next_state => N112, 
               clocked_on => CLK_port, Q => REGISTERS_43_28_port, QN => n_2379
               );
   REGISTERS_reg_43_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N135, next_state => N111, 
               clocked_on => CLK_port, Q => REGISTERS_43_27_port, QN => n_2380
               );
   REGISTERS_reg_43_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N135, next_state => N110, 
               clocked_on => CLK_port, Q => REGISTERS_43_26_port, QN => n_2381
               );
   REGISTERS_reg_43_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N135, next_state => N109, 
               clocked_on => CLK_port, Q => REGISTERS_43_25_port, QN => n_2382
               );
   REGISTERS_reg_43_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N135, next_state => N108, 
               clocked_on => CLK_port, Q => REGISTERS_43_24_port, QN => n_2383
               );
   REGISTERS_reg_43_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N135, next_state => N107, 
               clocked_on => CLK_port, Q => REGISTERS_43_23_port, QN => n_2384
               );
   REGISTERS_reg_43_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N135, next_state => N106, 
               clocked_on => CLK_port, Q => REGISTERS_43_22_port, QN => n_2385
               );
   REGISTERS_reg_43_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N135, next_state => N105, 
               clocked_on => CLK_port, Q => REGISTERS_43_21_port, QN => n_2386
               );
   REGISTERS_reg_43_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N135, next_state => N104, 
               clocked_on => CLK_port, Q => REGISTERS_43_20_port, QN => n_2387
               );
   REGISTERS_reg_43_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N135, next_state => N103, 
               clocked_on => CLK_port, Q => REGISTERS_43_19_port, QN => n_2388
               );
   REGISTERS_reg_43_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N135, next_state => N102, 
               clocked_on => CLK_port, Q => REGISTERS_43_18_port, QN => n_2389
               );
   REGISTERS_reg_43_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N135, next_state => N101, 
               clocked_on => CLK_port, Q => REGISTERS_43_17_port, QN => n_2390
               );
   REGISTERS_reg_43_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N135, next_state => N100, 
               clocked_on => CLK_port, Q => REGISTERS_43_16_port, QN => n_2391
               );
   REGISTERS_reg_43_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N135, next_state => N99, 
               clocked_on => CLK_port, Q => REGISTERS_43_15_port, QN => n_2392
               );
   REGISTERS_reg_43_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N135, next_state => N98, 
               clocked_on => CLK_port, Q => REGISTERS_43_14_port, QN => n_2393
               );
   REGISTERS_reg_43_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N135, next_state => N97, 
               clocked_on => CLK_port, Q => REGISTERS_43_13_port, QN => n_2394
               );
   REGISTERS_reg_43_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N135, next_state => N96, 
               clocked_on => CLK_port, Q => REGISTERS_43_12_port, QN => n_2395
               );
   REGISTERS_reg_43_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N135, next_state => N95, 
               clocked_on => CLK_port, Q => REGISTERS_43_11_port, QN => n_2396
               );
   REGISTERS_reg_43_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N135, next_state => N94, 
               clocked_on => CLK_port, Q => REGISTERS_43_10_port, QN => n_2397
               );
   REGISTERS_reg_43_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N135, next_state => N93, 
               clocked_on => CLK_port, Q => REGISTERS_43_9_port, QN => n_2398);
   REGISTERS_reg_43_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N135, next_state => N92, 
               clocked_on => CLK_port, Q => REGISTERS_43_8_port, QN => n_2399);
   REGISTERS_reg_43_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N135, next_state => N91, 
               clocked_on => CLK_port, Q => REGISTERS_43_7_port, QN => n_2400);
   REGISTERS_reg_43_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N135, next_state => N90, 
               clocked_on => CLK_port, Q => REGISTERS_43_6_port, QN => n_2401);
   REGISTERS_reg_43_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N135, next_state => N89, 
               clocked_on => CLK_port, Q => REGISTERS_43_5_port, QN => n_2402);
   REGISTERS_reg_43_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N135, next_state => N88, 
               clocked_on => CLK_port, Q => REGISTERS_43_4_port, QN => n_2403);
   REGISTERS_reg_43_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N135, next_state => N87, 
               clocked_on => CLK_port, Q => REGISTERS_43_3_port, QN => n_2404);
   REGISTERS_reg_43_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N135, next_state => N86, 
               clocked_on => CLK_port, Q => REGISTERS_43_2_port, QN => n_2405);
   REGISTERS_reg_43_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N135, next_state => N85, 
               clocked_on => CLK_port, Q => REGISTERS_43_1_port, QN => n_2406);
   REGISTERS_reg_43_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N135, next_state => N84, 
               clocked_on => CLK_port, Q => REGISTERS_43_0_port, QN => n_2407);
   REGISTERS_reg_44_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N134, next_state => N115, 
               clocked_on => CLK_port, Q => REGISTERS_44_31_port, QN => n_2408
               );
   REGISTERS_reg_44_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N134, next_state => N114, 
               clocked_on => CLK_port, Q => REGISTERS_44_30_port, QN => n_2409
               );
   REGISTERS_reg_44_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N134, next_state => N113, 
               clocked_on => CLK_port, Q => REGISTERS_44_29_port, QN => n_2410
               );
   REGISTERS_reg_44_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N134, next_state => N112, 
               clocked_on => CLK_port, Q => REGISTERS_44_28_port, QN => n_2411
               );
   REGISTERS_reg_44_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N134, next_state => N111, 
               clocked_on => CLK_port, Q => REGISTERS_44_27_port, QN => n_2412
               );
   REGISTERS_reg_44_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N134, next_state => N110, 
               clocked_on => CLK_port, Q => REGISTERS_44_26_port, QN => n_2413
               );
   REGISTERS_reg_44_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N134, next_state => N109, 
               clocked_on => CLK_port, Q => REGISTERS_44_25_port, QN => n_2414
               );
   REGISTERS_reg_44_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N134, next_state => N108, 
               clocked_on => CLK_port, Q => REGISTERS_44_24_port, QN => n_2415
               );
   REGISTERS_reg_44_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N134, next_state => N107, 
               clocked_on => CLK_port, Q => REGISTERS_44_23_port, QN => n_2416
               );
   REGISTERS_reg_44_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N134, next_state => N106, 
               clocked_on => CLK_port, Q => REGISTERS_44_22_port, QN => n_2417
               );
   REGISTERS_reg_44_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N134, next_state => N105, 
               clocked_on => CLK_port, Q => REGISTERS_44_21_port, QN => n_2418
               );
   REGISTERS_reg_44_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N134, next_state => N104, 
               clocked_on => CLK_port, Q => REGISTERS_44_20_port, QN => n_2419
               );
   REGISTERS_reg_44_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N134, next_state => N103, 
               clocked_on => CLK_port, Q => REGISTERS_44_19_port, QN => n_2420
               );
   REGISTERS_reg_44_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N134, next_state => N102, 
               clocked_on => CLK_port, Q => REGISTERS_44_18_port, QN => n_2421
               );
   REGISTERS_reg_44_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N134, next_state => N101, 
               clocked_on => CLK_port, Q => REGISTERS_44_17_port, QN => n_2422
               );
   REGISTERS_reg_44_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N134, next_state => N100, 
               clocked_on => CLK_port, Q => REGISTERS_44_16_port, QN => n_2423
               );
   REGISTERS_reg_44_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N134, next_state => N99, 
               clocked_on => CLK_port, Q => REGISTERS_44_15_port, QN => n_2424
               );
   REGISTERS_reg_44_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N134, next_state => N98, 
               clocked_on => CLK_port, Q => REGISTERS_44_14_port, QN => n_2425
               );
   REGISTERS_reg_44_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N134, next_state => N97, 
               clocked_on => CLK_port, Q => REGISTERS_44_13_port, QN => n_2426
               );
   REGISTERS_reg_44_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N134, next_state => N96, 
               clocked_on => CLK_port, Q => REGISTERS_44_12_port, QN => n_2427
               );
   REGISTERS_reg_44_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N134, next_state => N95, 
               clocked_on => CLK_port, Q => REGISTERS_44_11_port, QN => n_2428
               );
   REGISTERS_reg_44_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N134, next_state => N94, 
               clocked_on => CLK_port, Q => REGISTERS_44_10_port, QN => n_2429
               );
   REGISTERS_reg_44_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N134, next_state => N93, 
               clocked_on => CLK_port, Q => REGISTERS_44_9_port, QN => n_2430);
   REGISTERS_reg_44_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N134, next_state => N92, 
               clocked_on => CLK_port, Q => REGISTERS_44_8_port, QN => n_2431);
   REGISTERS_reg_44_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N134, next_state => N91, 
               clocked_on => CLK_port, Q => REGISTERS_44_7_port, QN => n_2432);
   REGISTERS_reg_44_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N134, next_state => N90, 
               clocked_on => CLK_port, Q => REGISTERS_44_6_port, QN => n_2433);
   REGISTERS_reg_44_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N134, next_state => N89, 
               clocked_on => CLK_port, Q => REGISTERS_44_5_port, QN => n_2434);
   REGISTERS_reg_44_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N134, next_state => N88, 
               clocked_on => CLK_port, Q => REGISTERS_44_4_port, QN => n_2435);
   REGISTERS_reg_44_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N134, next_state => N87, 
               clocked_on => CLK_port, Q => REGISTERS_44_3_port, QN => n_2436);
   REGISTERS_reg_44_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N134, next_state => N86, 
               clocked_on => CLK_port, Q => REGISTERS_44_2_port, QN => n_2437);
   REGISTERS_reg_44_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N134, next_state => N85, 
               clocked_on => CLK_port, Q => REGISTERS_44_1_port, QN => n_2438);
   REGISTERS_reg_44_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N134, next_state => N84, 
               clocked_on => CLK_port, Q => REGISTERS_44_0_port, QN => n_2439);
   REGISTERS_reg_45_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N133, next_state => N115, 
               clocked_on => CLK_port, Q => REGISTERS_45_31_port, QN => n_2440
               );
   REGISTERS_reg_45_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N133, next_state => N114, 
               clocked_on => CLK_port, Q => REGISTERS_45_30_port, QN => n_2441
               );
   REGISTERS_reg_45_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N133, next_state => N113, 
               clocked_on => CLK_port, Q => REGISTERS_45_29_port, QN => n_2442
               );
   REGISTERS_reg_45_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N133, next_state => N112, 
               clocked_on => CLK_port, Q => REGISTERS_45_28_port, QN => n_2443
               );
   REGISTERS_reg_45_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N133, next_state => N111, 
               clocked_on => CLK_port, Q => REGISTERS_45_27_port, QN => n_2444
               );
   REGISTERS_reg_45_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N133, next_state => N110, 
               clocked_on => CLK_port, Q => REGISTERS_45_26_port, QN => n_2445
               );
   REGISTERS_reg_45_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N133, next_state => N109, 
               clocked_on => CLK_port, Q => REGISTERS_45_25_port, QN => n_2446
               );
   REGISTERS_reg_45_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N133, next_state => N108, 
               clocked_on => CLK_port, Q => REGISTERS_45_24_port, QN => n_2447
               );
   REGISTERS_reg_45_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N133, next_state => N107, 
               clocked_on => CLK_port, Q => REGISTERS_45_23_port, QN => n_2448
               );
   REGISTERS_reg_45_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N133, next_state => N106, 
               clocked_on => CLK_port, Q => REGISTERS_45_22_port, QN => n_2449
               );
   REGISTERS_reg_45_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N133, next_state => N105, 
               clocked_on => CLK_port, Q => REGISTERS_45_21_port, QN => n_2450
               );
   REGISTERS_reg_45_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N133, next_state => N104, 
               clocked_on => CLK_port, Q => REGISTERS_45_20_port, QN => n_2451
               );
   REGISTERS_reg_45_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N133, next_state => N103, 
               clocked_on => CLK_port, Q => REGISTERS_45_19_port, QN => n_2452
               );
   REGISTERS_reg_45_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N133, next_state => N102, 
               clocked_on => CLK_port, Q => REGISTERS_45_18_port, QN => n_2453
               );
   REGISTERS_reg_45_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N133, next_state => N101, 
               clocked_on => CLK_port, Q => REGISTERS_45_17_port, QN => n_2454
               );
   REGISTERS_reg_45_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N133, next_state => N100, 
               clocked_on => CLK_port, Q => REGISTERS_45_16_port, QN => n_2455
               );
   REGISTERS_reg_45_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N133, next_state => N99, 
               clocked_on => CLK_port, Q => REGISTERS_45_15_port, QN => n_2456
               );
   REGISTERS_reg_45_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N133, next_state => N98, 
               clocked_on => CLK_port, Q => REGISTERS_45_14_port, QN => n_2457
               );
   REGISTERS_reg_45_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N133, next_state => N97, 
               clocked_on => CLK_port, Q => REGISTERS_45_13_port, QN => n_2458
               );
   REGISTERS_reg_45_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N133, next_state => N96, 
               clocked_on => CLK_port, Q => REGISTERS_45_12_port, QN => n_2459
               );
   REGISTERS_reg_45_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N133, next_state => N95, 
               clocked_on => CLK_port, Q => REGISTERS_45_11_port, QN => n_2460
               );
   REGISTERS_reg_45_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N133, next_state => N94, 
               clocked_on => CLK_port, Q => REGISTERS_45_10_port, QN => n_2461
               );
   REGISTERS_reg_45_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N133, next_state => N93, 
               clocked_on => CLK_port, Q => REGISTERS_45_9_port, QN => n_2462);
   REGISTERS_reg_45_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N133, next_state => N92, 
               clocked_on => CLK_port, Q => REGISTERS_45_8_port, QN => n_2463);
   REGISTERS_reg_45_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N133, next_state => N91, 
               clocked_on => CLK_port, Q => REGISTERS_45_7_port, QN => n_2464);
   REGISTERS_reg_45_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N133, next_state => N90, 
               clocked_on => CLK_port, Q => REGISTERS_45_6_port, QN => n_2465);
   REGISTERS_reg_45_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N133, next_state => N89, 
               clocked_on => CLK_port, Q => REGISTERS_45_5_port, QN => n_2466);
   REGISTERS_reg_45_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N133, next_state => N88, 
               clocked_on => CLK_port, Q => REGISTERS_45_4_port, QN => n_2467);
   REGISTERS_reg_45_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N133, next_state => N87, 
               clocked_on => CLK_port, Q => REGISTERS_45_3_port, QN => n_2468);
   REGISTERS_reg_45_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N133, next_state => N86, 
               clocked_on => CLK_port, Q => REGISTERS_45_2_port, QN => n_2469);
   REGISTERS_reg_45_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N133, next_state => N85, 
               clocked_on => CLK_port, Q => REGISTERS_45_1_port, QN => n_2470);
   REGISTERS_reg_45_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N133, next_state => N84, 
               clocked_on => CLK_port, Q => REGISTERS_45_0_port, QN => n_2471);
   REGISTERS_reg_46_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N132, next_state => N115, 
               clocked_on => CLK_port, Q => REGISTERS_46_31_port, QN => n_2472
               );
   REGISTERS_reg_46_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N132, next_state => N114, 
               clocked_on => CLK_port, Q => REGISTERS_46_30_port, QN => n_2473
               );
   REGISTERS_reg_46_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N132, next_state => N113, 
               clocked_on => CLK_port, Q => REGISTERS_46_29_port, QN => n_2474
               );
   REGISTERS_reg_46_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N132, next_state => N112, 
               clocked_on => CLK_port, Q => REGISTERS_46_28_port, QN => n_2475
               );
   REGISTERS_reg_46_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N132, next_state => N111, 
               clocked_on => CLK_port, Q => REGISTERS_46_27_port, QN => n_2476
               );
   REGISTERS_reg_46_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N132, next_state => N110, 
               clocked_on => CLK_port, Q => REGISTERS_46_26_port, QN => n_2477
               );
   REGISTERS_reg_46_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N132, next_state => N109, 
               clocked_on => CLK_port, Q => REGISTERS_46_25_port, QN => n_2478
               );
   REGISTERS_reg_46_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N132, next_state => N108, 
               clocked_on => CLK_port, Q => REGISTERS_46_24_port, QN => n_2479
               );
   REGISTERS_reg_46_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N132, next_state => N107, 
               clocked_on => CLK_port, Q => REGISTERS_46_23_port, QN => n_2480
               );
   REGISTERS_reg_46_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N132, next_state => N106, 
               clocked_on => CLK_port, Q => REGISTERS_46_22_port, QN => n_2481
               );
   REGISTERS_reg_46_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N132, next_state => N105, 
               clocked_on => CLK_port, Q => REGISTERS_46_21_port, QN => n_2482
               );
   REGISTERS_reg_46_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N132, next_state => N104, 
               clocked_on => CLK_port, Q => REGISTERS_46_20_port, QN => n_2483
               );
   REGISTERS_reg_46_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N132, next_state => N103, 
               clocked_on => CLK_port, Q => REGISTERS_46_19_port, QN => n_2484
               );
   REGISTERS_reg_46_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N132, next_state => N102, 
               clocked_on => CLK_port, Q => REGISTERS_46_18_port, QN => n_2485
               );
   REGISTERS_reg_46_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N132, next_state => N101, 
               clocked_on => CLK_port, Q => REGISTERS_46_17_port, QN => n_2486
               );
   REGISTERS_reg_46_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N132, next_state => N100, 
               clocked_on => CLK_port, Q => REGISTERS_46_16_port, QN => n_2487
               );
   REGISTERS_reg_46_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N132, next_state => N99, 
               clocked_on => CLK_port, Q => REGISTERS_46_15_port, QN => n_2488
               );
   REGISTERS_reg_46_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N132, next_state => N98, 
               clocked_on => CLK_port, Q => REGISTERS_46_14_port, QN => n_2489
               );
   REGISTERS_reg_46_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N132, next_state => N97, 
               clocked_on => CLK_port, Q => REGISTERS_46_13_port, QN => n_2490
               );
   REGISTERS_reg_46_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N132, next_state => N96, 
               clocked_on => CLK_port, Q => REGISTERS_46_12_port, QN => n_2491
               );
   REGISTERS_reg_46_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N132, next_state => N95, 
               clocked_on => CLK_port, Q => REGISTERS_46_11_port, QN => n_2492
               );
   REGISTERS_reg_46_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N132, next_state => N94, 
               clocked_on => CLK_port, Q => REGISTERS_46_10_port, QN => n_2493
               );
   REGISTERS_reg_46_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N132, next_state => N93, 
               clocked_on => CLK_port, Q => REGISTERS_46_9_port, QN => n_2494);
   REGISTERS_reg_46_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N132, next_state => N92, 
               clocked_on => CLK_port, Q => REGISTERS_46_8_port, QN => n_2495);
   REGISTERS_reg_46_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N132, next_state => N91, 
               clocked_on => CLK_port, Q => REGISTERS_46_7_port, QN => n_2496);
   REGISTERS_reg_46_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N132, next_state => N90, 
               clocked_on => CLK_port, Q => REGISTERS_46_6_port, QN => n_2497);
   REGISTERS_reg_46_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N132, next_state => N89, 
               clocked_on => CLK_port, Q => REGISTERS_46_5_port, QN => n_2498);
   REGISTERS_reg_46_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N132, next_state => N88, 
               clocked_on => CLK_port, Q => REGISTERS_46_4_port, QN => n_2499);
   REGISTERS_reg_46_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N132, next_state => N87, 
               clocked_on => CLK_port, Q => REGISTERS_46_3_port, QN => n_2500);
   REGISTERS_reg_46_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N132, next_state => N86, 
               clocked_on => CLK_port, Q => REGISTERS_46_2_port, QN => n_2501);
   REGISTERS_reg_46_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N132, next_state => N85, 
               clocked_on => CLK_port, Q => REGISTERS_46_1_port, QN => n_2502);
   REGISTERS_reg_46_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N132, next_state => N84, 
               clocked_on => CLK_port, Q => REGISTERS_46_0_port, QN => n_2503);
   REGISTERS_reg_47_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N131, next_state => N115, 
               clocked_on => CLK_port, Q => REGISTERS_47_31_port, QN => n_2504
               );
   REGISTERS_reg_47_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N131, next_state => N114, 
               clocked_on => CLK_port, Q => REGISTERS_47_30_port, QN => n_2505
               );
   REGISTERS_reg_47_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N131, next_state => N113, 
               clocked_on => CLK_port, Q => REGISTERS_47_29_port, QN => n_2506
               );
   REGISTERS_reg_47_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N131, next_state => N112, 
               clocked_on => CLK_port, Q => REGISTERS_47_28_port, QN => n_2507
               );
   REGISTERS_reg_47_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N131, next_state => N111, 
               clocked_on => CLK_port, Q => REGISTERS_47_27_port, QN => n_2508
               );
   REGISTERS_reg_47_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N131, next_state => N110, 
               clocked_on => CLK_port, Q => REGISTERS_47_26_port, QN => n_2509
               );
   REGISTERS_reg_47_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N131, next_state => N109, 
               clocked_on => CLK_port, Q => REGISTERS_47_25_port, QN => n_2510
               );
   REGISTERS_reg_47_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N131, next_state => N108, 
               clocked_on => CLK_port, Q => REGISTERS_47_24_port, QN => n_2511
               );
   REGISTERS_reg_47_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N131, next_state => N107, 
               clocked_on => CLK_port, Q => REGISTERS_47_23_port, QN => n_2512
               );
   REGISTERS_reg_47_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N131, next_state => N106, 
               clocked_on => CLK_port, Q => REGISTERS_47_22_port, QN => n_2513
               );
   REGISTERS_reg_47_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N131, next_state => N105, 
               clocked_on => CLK_port, Q => REGISTERS_47_21_port, QN => n_2514
               );
   REGISTERS_reg_47_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N131, next_state => N104, 
               clocked_on => CLK_port, Q => REGISTERS_47_20_port, QN => n_2515
               );
   REGISTERS_reg_47_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N131, next_state => N103, 
               clocked_on => CLK_port, Q => REGISTERS_47_19_port, QN => n_2516
               );
   REGISTERS_reg_47_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N131, next_state => N102, 
               clocked_on => CLK_port, Q => REGISTERS_47_18_port, QN => n_2517
               );
   REGISTERS_reg_47_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N131, next_state => N101, 
               clocked_on => CLK_port, Q => REGISTERS_47_17_port, QN => n_2518
               );
   REGISTERS_reg_47_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N131, next_state => N100, 
               clocked_on => CLK_port, Q => REGISTERS_47_16_port, QN => n_2519
               );
   REGISTERS_reg_47_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N131, next_state => N99, 
               clocked_on => CLK_port, Q => REGISTERS_47_15_port, QN => n_2520
               );
   REGISTERS_reg_47_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N131, next_state => N98, 
               clocked_on => CLK_port, Q => REGISTERS_47_14_port, QN => n_2521
               );
   REGISTERS_reg_47_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N131, next_state => N97, 
               clocked_on => CLK_port, Q => REGISTERS_47_13_port, QN => n_2522
               );
   REGISTERS_reg_47_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N131, next_state => N96, 
               clocked_on => CLK_port, Q => REGISTERS_47_12_port, QN => n_2523
               );
   REGISTERS_reg_47_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N131, next_state => N95, 
               clocked_on => CLK_port, Q => REGISTERS_47_11_port, QN => n_2524
               );
   REGISTERS_reg_47_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N131, next_state => N94, 
               clocked_on => CLK_port, Q => REGISTERS_47_10_port, QN => n_2525
               );
   REGISTERS_reg_47_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N131, next_state => N93, 
               clocked_on => CLK_port, Q => REGISTERS_47_9_port, QN => n_2526);
   REGISTERS_reg_47_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N131, next_state => N92, 
               clocked_on => CLK_port, Q => REGISTERS_47_8_port, QN => n_2527);
   REGISTERS_reg_47_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N131, next_state => N91, 
               clocked_on => CLK_port, Q => REGISTERS_47_7_port, QN => n_2528);
   REGISTERS_reg_47_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N131, next_state => N90, 
               clocked_on => CLK_port, Q => REGISTERS_47_6_port, QN => n_2529);
   REGISTERS_reg_47_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N131, next_state => N89, 
               clocked_on => CLK_port, Q => REGISTERS_47_5_port, QN => n_2530);
   REGISTERS_reg_47_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N131, next_state => N88, 
               clocked_on => CLK_port, Q => REGISTERS_47_4_port, QN => n_2531);
   REGISTERS_reg_47_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N131, next_state => N87, 
               clocked_on => CLK_port, Q => REGISTERS_47_3_port, QN => n_2532);
   REGISTERS_reg_47_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N131, next_state => N86, 
               clocked_on => CLK_port, Q => REGISTERS_47_2_port, QN => n_2533);
   REGISTERS_reg_47_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N131, next_state => N85, 
               clocked_on => CLK_port, Q => REGISTERS_47_1_port, QN => n_2534);
   REGISTERS_reg_47_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N131, next_state => N84, 
               clocked_on => CLK_port, Q => REGISTERS_47_0_port, QN => n_2535);
   REGISTERS_reg_48_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N130, next_state => N115, 
               clocked_on => CLK_port, Q => REGISTERS_48_31_port, QN => n_2536
               );
   REGISTERS_reg_48_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N130, next_state => N114, 
               clocked_on => CLK_port, Q => REGISTERS_48_30_port, QN => n_2537
               );
   REGISTERS_reg_48_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N130, next_state => N113, 
               clocked_on => CLK_port, Q => REGISTERS_48_29_port, QN => n_2538
               );
   REGISTERS_reg_48_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N130, next_state => N112, 
               clocked_on => CLK_port, Q => REGISTERS_48_28_port, QN => n_2539
               );
   REGISTERS_reg_48_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N130, next_state => N111, 
               clocked_on => CLK_port, Q => REGISTERS_48_27_port, QN => n_2540
               );
   REGISTERS_reg_48_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N130, next_state => N110, 
               clocked_on => CLK_port, Q => REGISTERS_48_26_port, QN => n_2541
               );
   REGISTERS_reg_48_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N130, next_state => N109, 
               clocked_on => CLK_port, Q => REGISTERS_48_25_port, QN => n_2542
               );
   REGISTERS_reg_48_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N130, next_state => N108, 
               clocked_on => CLK_port, Q => REGISTERS_48_24_port, QN => n_2543
               );
   REGISTERS_reg_48_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N130, next_state => N107, 
               clocked_on => CLK_port, Q => REGISTERS_48_23_port, QN => n_2544
               );
   REGISTERS_reg_48_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N130, next_state => N106, 
               clocked_on => CLK_port, Q => REGISTERS_48_22_port, QN => n_2545
               );
   REGISTERS_reg_48_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N130, next_state => N105, 
               clocked_on => CLK_port, Q => REGISTERS_48_21_port, QN => n_2546
               );
   REGISTERS_reg_48_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N130, next_state => N104, 
               clocked_on => CLK_port, Q => REGISTERS_48_20_port, QN => n_2547
               );
   REGISTERS_reg_48_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N130, next_state => N103, 
               clocked_on => CLK_port, Q => REGISTERS_48_19_port, QN => n_2548
               );
   REGISTERS_reg_48_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N130, next_state => N102, 
               clocked_on => CLK_port, Q => REGISTERS_48_18_port, QN => n_2549
               );
   REGISTERS_reg_48_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N130, next_state => N101, 
               clocked_on => CLK_port, Q => REGISTERS_48_17_port, QN => n_2550
               );
   REGISTERS_reg_48_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N130, next_state => N100, 
               clocked_on => CLK_port, Q => REGISTERS_48_16_port, QN => n_2551
               );
   REGISTERS_reg_48_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N130, next_state => N99, 
               clocked_on => CLK_port, Q => REGISTERS_48_15_port, QN => n_2552
               );
   REGISTERS_reg_48_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N130, next_state => N98, 
               clocked_on => CLK_port, Q => REGISTERS_48_14_port, QN => n_2553
               );
   REGISTERS_reg_48_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N130, next_state => N97, 
               clocked_on => CLK_port, Q => REGISTERS_48_13_port, QN => n_2554
               );
   REGISTERS_reg_48_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N130, next_state => N96, 
               clocked_on => CLK_port, Q => REGISTERS_48_12_port, QN => n_2555
               );
   REGISTERS_reg_48_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N130, next_state => N95, 
               clocked_on => CLK_port, Q => REGISTERS_48_11_port, QN => n_2556
               );
   REGISTERS_reg_48_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N130, next_state => N94, 
               clocked_on => CLK_port, Q => REGISTERS_48_10_port, QN => n_2557
               );
   REGISTERS_reg_48_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N130, next_state => N93, 
               clocked_on => CLK_port, Q => REGISTERS_48_9_port, QN => n_2558);
   REGISTERS_reg_48_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N130, next_state => N92, 
               clocked_on => CLK_port, Q => REGISTERS_48_8_port, QN => n_2559);
   REGISTERS_reg_48_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N130, next_state => N91, 
               clocked_on => CLK_port, Q => REGISTERS_48_7_port, QN => n_2560);
   REGISTERS_reg_48_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N130, next_state => N90, 
               clocked_on => CLK_port, Q => REGISTERS_48_6_port, QN => n_2561);
   REGISTERS_reg_48_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N130, next_state => N89, 
               clocked_on => CLK_port, Q => REGISTERS_48_5_port, QN => n_2562);
   REGISTERS_reg_48_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N130, next_state => N88, 
               clocked_on => CLK_port, Q => REGISTERS_48_4_port, QN => n_2563);
   REGISTERS_reg_48_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N130, next_state => N87, 
               clocked_on => CLK_port, Q => REGISTERS_48_3_port, QN => n_2564);
   REGISTERS_reg_48_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N130, next_state => N86, 
               clocked_on => CLK_port, Q => REGISTERS_48_2_port, QN => n_2565);
   REGISTERS_reg_48_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N130, next_state => N85, 
               clocked_on => CLK_port, Q => REGISTERS_48_1_port, QN => n_2566);
   REGISTERS_reg_48_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N130, next_state => N84, 
               clocked_on => CLK_port, Q => REGISTERS_48_0_port, QN => n_2567);
   REGISTERS_reg_49_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N129, next_state => N115, 
               clocked_on => CLK_port, Q => REGISTERS_49_31_port, QN => n_2568
               );
   REGISTERS_reg_49_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N129, next_state => N114, 
               clocked_on => CLK_port, Q => REGISTERS_49_30_port, QN => n_2569
               );
   REGISTERS_reg_49_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N129, next_state => N113, 
               clocked_on => CLK_port, Q => REGISTERS_49_29_port, QN => n_2570
               );
   REGISTERS_reg_49_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N129, next_state => N112, 
               clocked_on => CLK_port, Q => REGISTERS_49_28_port, QN => n_2571
               );
   REGISTERS_reg_49_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N129, next_state => N111, 
               clocked_on => CLK_port, Q => REGISTERS_49_27_port, QN => n_2572
               );
   REGISTERS_reg_49_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N129, next_state => N110, 
               clocked_on => CLK_port, Q => REGISTERS_49_26_port, QN => n_2573
               );
   REGISTERS_reg_49_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N129, next_state => N109, 
               clocked_on => CLK_port, Q => REGISTERS_49_25_port, QN => n_2574
               );
   REGISTERS_reg_49_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N129, next_state => N108, 
               clocked_on => CLK_port, Q => REGISTERS_49_24_port, QN => n_2575
               );
   REGISTERS_reg_49_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N129, next_state => N107, 
               clocked_on => CLK_port, Q => REGISTERS_49_23_port, QN => n_2576
               );
   REGISTERS_reg_49_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N129, next_state => N106, 
               clocked_on => CLK_port, Q => REGISTERS_49_22_port, QN => n_2577
               );
   REGISTERS_reg_49_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N129, next_state => N105, 
               clocked_on => CLK_port, Q => REGISTERS_49_21_port, QN => n_2578
               );
   REGISTERS_reg_49_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N129, next_state => N104, 
               clocked_on => CLK_port, Q => REGISTERS_49_20_port, QN => n_2579
               );
   REGISTERS_reg_49_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N129, next_state => N103, 
               clocked_on => CLK_port, Q => REGISTERS_49_19_port, QN => n_2580
               );
   REGISTERS_reg_49_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N129, next_state => N102, 
               clocked_on => CLK_port, Q => REGISTERS_49_18_port, QN => n_2581
               );
   REGISTERS_reg_49_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N129, next_state => N101, 
               clocked_on => CLK_port, Q => REGISTERS_49_17_port, QN => n_2582
               );
   REGISTERS_reg_49_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N129, next_state => N100, 
               clocked_on => CLK_port, Q => REGISTERS_49_16_port, QN => n_2583
               );
   REGISTERS_reg_49_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N129, next_state => N99, 
               clocked_on => CLK_port, Q => REGISTERS_49_15_port, QN => n_2584
               );
   REGISTERS_reg_49_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N129, next_state => N98, 
               clocked_on => CLK_port, Q => REGISTERS_49_14_port, QN => n_2585
               );
   REGISTERS_reg_49_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N129, next_state => N97, 
               clocked_on => CLK_port, Q => REGISTERS_49_13_port, QN => n_2586
               );
   REGISTERS_reg_49_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N129, next_state => N96, 
               clocked_on => CLK_port, Q => REGISTERS_49_12_port, QN => n_2587
               );
   REGISTERS_reg_49_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N129, next_state => N95, 
               clocked_on => CLK_port, Q => REGISTERS_49_11_port, QN => n_2588
               );
   REGISTERS_reg_49_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N129, next_state => N94, 
               clocked_on => CLK_port, Q => REGISTERS_49_10_port, QN => n_2589
               );
   REGISTERS_reg_49_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N129, next_state => N93, 
               clocked_on => CLK_port, Q => REGISTERS_49_9_port, QN => n_2590);
   REGISTERS_reg_49_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N129, next_state => N92, 
               clocked_on => CLK_port, Q => REGISTERS_49_8_port, QN => n_2591);
   REGISTERS_reg_49_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N129, next_state => N91, 
               clocked_on => CLK_port, Q => REGISTERS_49_7_port, QN => n_2592);
   REGISTERS_reg_49_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N129, next_state => N90, 
               clocked_on => CLK_port, Q => REGISTERS_49_6_port, QN => n_2593);
   REGISTERS_reg_49_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N129, next_state => N89, 
               clocked_on => CLK_port, Q => REGISTERS_49_5_port, QN => n_2594);
   REGISTERS_reg_49_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N129, next_state => N88, 
               clocked_on => CLK_port, Q => REGISTERS_49_4_port, QN => n_2595);
   REGISTERS_reg_49_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N129, next_state => N87, 
               clocked_on => CLK_port, Q => REGISTERS_49_3_port, QN => n_2596);
   REGISTERS_reg_49_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N129, next_state => N86, 
               clocked_on => CLK_port, Q => REGISTERS_49_2_port, QN => n_2597);
   REGISTERS_reg_49_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N129, next_state => N85, 
               clocked_on => CLK_port, Q => REGISTERS_49_1_port, QN => n_2598);
   REGISTERS_reg_49_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N129, next_state => N84, 
               clocked_on => CLK_port, Q => REGISTERS_49_0_port, QN => n_2599);
   REGISTERS_reg_50_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N128, next_state => N115, 
               clocked_on => CLK_port, Q => REGISTERS_50_31_port, QN => n_2600
               );
   REGISTERS_reg_50_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N128, next_state => N114, 
               clocked_on => CLK_port, Q => REGISTERS_50_30_port, QN => n_2601
               );
   REGISTERS_reg_50_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N128, next_state => N113, 
               clocked_on => CLK_port, Q => REGISTERS_50_29_port, QN => n_2602
               );
   REGISTERS_reg_50_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N128, next_state => N112, 
               clocked_on => CLK_port, Q => REGISTERS_50_28_port, QN => n_2603
               );
   REGISTERS_reg_50_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N128, next_state => N111, 
               clocked_on => CLK_port, Q => REGISTERS_50_27_port, QN => n_2604
               );
   REGISTERS_reg_50_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N128, next_state => N110, 
               clocked_on => CLK_port, Q => REGISTERS_50_26_port, QN => n_2605
               );
   REGISTERS_reg_50_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N128, next_state => N109, 
               clocked_on => CLK_port, Q => REGISTERS_50_25_port, QN => n_2606
               );
   REGISTERS_reg_50_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N128, next_state => N108, 
               clocked_on => CLK_port, Q => REGISTERS_50_24_port, QN => n_2607
               );
   REGISTERS_reg_50_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N128, next_state => N107, 
               clocked_on => CLK_port, Q => REGISTERS_50_23_port, QN => n_2608
               );
   REGISTERS_reg_50_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N128, next_state => N106, 
               clocked_on => CLK_port, Q => REGISTERS_50_22_port, QN => n_2609
               );
   REGISTERS_reg_50_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N128, next_state => N105, 
               clocked_on => CLK_port, Q => REGISTERS_50_21_port, QN => n_2610
               );
   REGISTERS_reg_50_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N128, next_state => N104, 
               clocked_on => CLK_port, Q => REGISTERS_50_20_port, QN => n_2611
               );
   REGISTERS_reg_50_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N128, next_state => N103, 
               clocked_on => CLK_port, Q => REGISTERS_50_19_port, QN => n_2612
               );
   REGISTERS_reg_50_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N128, next_state => N102, 
               clocked_on => CLK_port, Q => REGISTERS_50_18_port, QN => n_2613
               );
   REGISTERS_reg_50_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N128, next_state => N101, 
               clocked_on => CLK_port, Q => REGISTERS_50_17_port, QN => n_2614
               );
   REGISTERS_reg_50_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N128, next_state => N100, 
               clocked_on => CLK_port, Q => REGISTERS_50_16_port, QN => n_2615
               );
   REGISTERS_reg_50_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N128, next_state => N99, 
               clocked_on => CLK_port, Q => REGISTERS_50_15_port, QN => n_2616
               );
   REGISTERS_reg_50_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N128, next_state => N98, 
               clocked_on => CLK_port, Q => REGISTERS_50_14_port, QN => n_2617
               );
   REGISTERS_reg_50_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N128, next_state => N97, 
               clocked_on => CLK_port, Q => REGISTERS_50_13_port, QN => n_2618
               );
   REGISTERS_reg_50_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N128, next_state => N96, 
               clocked_on => CLK_port, Q => REGISTERS_50_12_port, QN => n_2619
               );
   REGISTERS_reg_50_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N128, next_state => N95, 
               clocked_on => CLK_port, Q => REGISTERS_50_11_port, QN => n_2620
               );
   REGISTERS_reg_50_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N128, next_state => N94, 
               clocked_on => CLK_port, Q => REGISTERS_50_10_port, QN => n_2621
               );
   REGISTERS_reg_50_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N128, next_state => N93, 
               clocked_on => CLK_port, Q => REGISTERS_50_9_port, QN => n_2622);
   REGISTERS_reg_50_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N128, next_state => N92, 
               clocked_on => CLK_port, Q => REGISTERS_50_8_port, QN => n_2623);
   REGISTERS_reg_50_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N128, next_state => N91, 
               clocked_on => CLK_port, Q => REGISTERS_50_7_port, QN => n_2624);
   REGISTERS_reg_50_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N128, next_state => N90, 
               clocked_on => CLK_port, Q => REGISTERS_50_6_port, QN => n_2625);
   REGISTERS_reg_50_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N128, next_state => N89, 
               clocked_on => CLK_port, Q => REGISTERS_50_5_port, QN => n_2626);
   REGISTERS_reg_50_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N128, next_state => N88, 
               clocked_on => CLK_port, Q => REGISTERS_50_4_port, QN => n_2627);
   REGISTERS_reg_50_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N128, next_state => N87, 
               clocked_on => CLK_port, Q => REGISTERS_50_3_port, QN => n_2628);
   REGISTERS_reg_50_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N128, next_state => N86, 
               clocked_on => CLK_port, Q => REGISTERS_50_2_port, QN => n_2629);
   REGISTERS_reg_50_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N128, next_state => N85, 
               clocked_on => CLK_port, Q => REGISTERS_50_1_port, QN => n_2630);
   REGISTERS_reg_50_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N128, next_state => N84, 
               clocked_on => CLK_port, Q => REGISTERS_50_0_port, QN => n_2631);
   REGISTERS_reg_51_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N127, next_state => N115, 
               clocked_on => CLK_port, Q => REGISTERS_51_31_port, QN => n_2632
               );
   REGISTERS_reg_51_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N127, next_state => N114, 
               clocked_on => CLK_port, Q => REGISTERS_51_30_port, QN => n_2633
               );
   REGISTERS_reg_51_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N127, next_state => N113, 
               clocked_on => CLK_port, Q => REGISTERS_51_29_port, QN => n_2634
               );
   REGISTERS_reg_51_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N127, next_state => N112, 
               clocked_on => CLK_port, Q => REGISTERS_51_28_port, QN => n_2635
               );
   REGISTERS_reg_51_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N127, next_state => N111, 
               clocked_on => CLK_port, Q => REGISTERS_51_27_port, QN => n_2636
               );
   REGISTERS_reg_51_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N127, next_state => N110, 
               clocked_on => CLK_port, Q => REGISTERS_51_26_port, QN => n_2637
               );
   REGISTERS_reg_51_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N127, next_state => N109, 
               clocked_on => CLK_port, Q => REGISTERS_51_25_port, QN => n_2638
               );
   REGISTERS_reg_51_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N127, next_state => N108, 
               clocked_on => CLK_port, Q => REGISTERS_51_24_port, QN => n_2639
               );
   REGISTERS_reg_51_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N127, next_state => N107, 
               clocked_on => CLK_port, Q => REGISTERS_51_23_port, QN => n_2640
               );
   REGISTERS_reg_51_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N127, next_state => N106, 
               clocked_on => CLK_port, Q => REGISTERS_51_22_port, QN => n_2641
               );
   REGISTERS_reg_51_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N127, next_state => N105, 
               clocked_on => CLK_port, Q => REGISTERS_51_21_port, QN => n_2642
               );
   REGISTERS_reg_51_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N127, next_state => N104, 
               clocked_on => CLK_port, Q => REGISTERS_51_20_port, QN => n_2643
               );
   REGISTERS_reg_51_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N127, next_state => N103, 
               clocked_on => CLK_port, Q => REGISTERS_51_19_port, QN => n_2644
               );
   REGISTERS_reg_51_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N127, next_state => N102, 
               clocked_on => CLK_port, Q => REGISTERS_51_18_port, QN => n_2645
               );
   REGISTERS_reg_51_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N127, next_state => N101, 
               clocked_on => CLK_port, Q => REGISTERS_51_17_port, QN => n_2646
               );
   REGISTERS_reg_51_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N127, next_state => N100, 
               clocked_on => CLK_port, Q => REGISTERS_51_16_port, QN => n_2647
               );
   REGISTERS_reg_51_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N127, next_state => N99, 
               clocked_on => CLK_port, Q => REGISTERS_51_15_port, QN => n_2648
               );
   REGISTERS_reg_51_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N127, next_state => N98, 
               clocked_on => CLK_port, Q => REGISTERS_51_14_port, QN => n_2649
               );
   REGISTERS_reg_51_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N127, next_state => N97, 
               clocked_on => CLK_port, Q => REGISTERS_51_13_port, QN => n_2650
               );
   REGISTERS_reg_51_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N127, next_state => N96, 
               clocked_on => CLK_port, Q => REGISTERS_51_12_port, QN => n_2651
               );
   REGISTERS_reg_51_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N127, next_state => N95, 
               clocked_on => CLK_port, Q => REGISTERS_51_11_port, QN => n_2652
               );
   REGISTERS_reg_51_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N127, next_state => N94, 
               clocked_on => CLK_port, Q => REGISTERS_51_10_port, QN => n_2653
               );
   REGISTERS_reg_51_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N127, next_state => N93, 
               clocked_on => CLK_port, Q => REGISTERS_51_9_port, QN => n_2654);
   REGISTERS_reg_51_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N127, next_state => N92, 
               clocked_on => CLK_port, Q => REGISTERS_51_8_port, QN => n_2655);
   REGISTERS_reg_51_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N127, next_state => N91, 
               clocked_on => CLK_port, Q => REGISTERS_51_7_port, QN => n_2656);
   REGISTERS_reg_51_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N127, next_state => N90, 
               clocked_on => CLK_port, Q => REGISTERS_51_6_port, QN => n_2657);
   REGISTERS_reg_51_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N127, next_state => N89, 
               clocked_on => CLK_port, Q => REGISTERS_51_5_port, QN => n_2658);
   REGISTERS_reg_51_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N127, next_state => N88, 
               clocked_on => CLK_port, Q => REGISTERS_51_4_port, QN => n_2659);
   REGISTERS_reg_51_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N127, next_state => N87, 
               clocked_on => CLK_port, Q => REGISTERS_51_3_port, QN => n_2660);
   REGISTERS_reg_51_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N127, next_state => N86, 
               clocked_on => CLK_port, Q => REGISTERS_51_2_port, QN => n_2661);
   REGISTERS_reg_51_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N127, next_state => N85, 
               clocked_on => CLK_port, Q => REGISTERS_51_1_port, QN => n_2662);
   REGISTERS_reg_51_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N127, next_state => N84, 
               clocked_on => CLK_port, Q => REGISTERS_51_0_port, QN => n_2663);
   REGISTERS_reg_52_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N126, next_state => N115, 
               clocked_on => CLK_port, Q => REGISTERS_52_31_port, QN => n_2664
               );
   REGISTERS_reg_52_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N126, next_state => N114, 
               clocked_on => CLK_port, Q => REGISTERS_52_30_port, QN => n_2665
               );
   REGISTERS_reg_52_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N126, next_state => N113, 
               clocked_on => CLK_port, Q => REGISTERS_52_29_port, QN => n_2666
               );
   REGISTERS_reg_52_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N126, next_state => N112, 
               clocked_on => CLK_port, Q => REGISTERS_52_28_port, QN => n_2667
               );
   REGISTERS_reg_52_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N126, next_state => N111, 
               clocked_on => CLK_port, Q => REGISTERS_52_27_port, QN => n_2668
               );
   REGISTERS_reg_52_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N126, next_state => N110, 
               clocked_on => CLK_port, Q => REGISTERS_52_26_port, QN => n_2669
               );
   REGISTERS_reg_52_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N126, next_state => N109, 
               clocked_on => CLK_port, Q => REGISTERS_52_25_port, QN => n_2670
               );
   REGISTERS_reg_52_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N126, next_state => N108, 
               clocked_on => CLK_port, Q => REGISTERS_52_24_port, QN => n_2671
               );
   REGISTERS_reg_52_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N126, next_state => N107, 
               clocked_on => CLK_port, Q => REGISTERS_52_23_port, QN => n_2672
               );
   REGISTERS_reg_52_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N126, next_state => N106, 
               clocked_on => CLK_port, Q => REGISTERS_52_22_port, QN => n_2673
               );
   REGISTERS_reg_52_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N126, next_state => N105, 
               clocked_on => CLK_port, Q => REGISTERS_52_21_port, QN => n_2674
               );
   REGISTERS_reg_52_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N126, next_state => N104, 
               clocked_on => CLK_port, Q => REGISTERS_52_20_port, QN => n_2675
               );
   REGISTERS_reg_52_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N126, next_state => N103, 
               clocked_on => CLK_port, Q => REGISTERS_52_19_port, QN => n_2676
               );
   REGISTERS_reg_52_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N126, next_state => N102, 
               clocked_on => CLK_port, Q => REGISTERS_52_18_port, QN => n_2677
               );
   REGISTERS_reg_52_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N126, next_state => N101, 
               clocked_on => CLK_port, Q => REGISTERS_52_17_port, QN => n_2678
               );
   REGISTERS_reg_52_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N126, next_state => N100, 
               clocked_on => CLK_port, Q => REGISTERS_52_16_port, QN => n_2679
               );
   REGISTERS_reg_52_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N126, next_state => N99, 
               clocked_on => CLK_port, Q => REGISTERS_52_15_port, QN => n_2680
               );
   REGISTERS_reg_52_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N126, next_state => N98, 
               clocked_on => CLK_port, Q => REGISTERS_52_14_port, QN => n_2681
               );
   REGISTERS_reg_52_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N126, next_state => N97, 
               clocked_on => CLK_port, Q => REGISTERS_52_13_port, QN => n_2682
               );
   REGISTERS_reg_52_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N126, next_state => N96, 
               clocked_on => CLK_port, Q => REGISTERS_52_12_port, QN => n_2683
               );
   REGISTERS_reg_52_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N126, next_state => N95, 
               clocked_on => CLK_port, Q => REGISTERS_52_11_port, QN => n_2684
               );
   REGISTERS_reg_52_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N126, next_state => N94, 
               clocked_on => CLK_port, Q => REGISTERS_52_10_port, QN => n_2685
               );
   REGISTERS_reg_52_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N126, next_state => N93, 
               clocked_on => CLK_port, Q => REGISTERS_52_9_port, QN => n_2686);
   REGISTERS_reg_52_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N126, next_state => N92, 
               clocked_on => CLK_port, Q => REGISTERS_52_8_port, QN => n_2687);
   REGISTERS_reg_52_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N126, next_state => N91, 
               clocked_on => CLK_port, Q => REGISTERS_52_7_port, QN => n_2688);
   REGISTERS_reg_52_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N126, next_state => N90, 
               clocked_on => CLK_port, Q => REGISTERS_52_6_port, QN => n_2689);
   REGISTERS_reg_52_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N126, next_state => N89, 
               clocked_on => CLK_port, Q => REGISTERS_52_5_port, QN => n_2690);
   REGISTERS_reg_52_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N126, next_state => N88, 
               clocked_on => CLK_port, Q => REGISTERS_52_4_port, QN => n_2691);
   REGISTERS_reg_52_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N126, next_state => N87, 
               clocked_on => CLK_port, Q => REGISTERS_52_3_port, QN => n_2692);
   REGISTERS_reg_52_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N126, next_state => N86, 
               clocked_on => CLK_port, Q => REGISTERS_52_2_port, QN => n_2693);
   REGISTERS_reg_52_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N126, next_state => N85, 
               clocked_on => CLK_port, Q => REGISTERS_52_1_port, QN => n_2694);
   REGISTERS_reg_52_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N126, next_state => N84, 
               clocked_on => CLK_port, Q => REGISTERS_52_0_port, QN => n_2695);
   REGISTERS_reg_53_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N125, next_state => N115, 
               clocked_on => CLK_port, Q => REGISTERS_53_31_port, QN => n_2696
               );
   REGISTERS_reg_53_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N125, next_state => N114, 
               clocked_on => CLK_port, Q => REGISTERS_53_30_port, QN => n_2697
               );
   REGISTERS_reg_53_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N125, next_state => N113, 
               clocked_on => CLK_port, Q => REGISTERS_53_29_port, QN => n_2698
               );
   REGISTERS_reg_53_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N125, next_state => N112, 
               clocked_on => CLK_port, Q => REGISTERS_53_28_port, QN => n_2699
               );
   REGISTERS_reg_53_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N125, next_state => N111, 
               clocked_on => CLK_port, Q => REGISTERS_53_27_port, QN => n_2700
               );
   REGISTERS_reg_53_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N125, next_state => N110, 
               clocked_on => CLK_port, Q => REGISTERS_53_26_port, QN => n_2701
               );
   REGISTERS_reg_53_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N125, next_state => N109, 
               clocked_on => CLK_port, Q => REGISTERS_53_25_port, QN => n_2702
               );
   REGISTERS_reg_53_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N125, next_state => N108, 
               clocked_on => CLK_port, Q => REGISTERS_53_24_port, QN => n_2703
               );
   REGISTERS_reg_53_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N125, next_state => N107, 
               clocked_on => CLK_port, Q => REGISTERS_53_23_port, QN => n_2704
               );
   REGISTERS_reg_53_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N125, next_state => N106, 
               clocked_on => CLK_port, Q => REGISTERS_53_22_port, QN => n_2705
               );
   REGISTERS_reg_53_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N125, next_state => N105, 
               clocked_on => CLK_port, Q => REGISTERS_53_21_port, QN => n_2706
               );
   REGISTERS_reg_53_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N125, next_state => N104, 
               clocked_on => CLK_port, Q => REGISTERS_53_20_port, QN => n_2707
               );
   REGISTERS_reg_53_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N125, next_state => N103, 
               clocked_on => CLK_port, Q => REGISTERS_53_19_port, QN => n_2708
               );
   REGISTERS_reg_53_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N125, next_state => N102, 
               clocked_on => CLK_port, Q => REGISTERS_53_18_port, QN => n_2709
               );
   REGISTERS_reg_53_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N125, next_state => N101, 
               clocked_on => CLK_port, Q => REGISTERS_53_17_port, QN => n_2710
               );
   REGISTERS_reg_53_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N125, next_state => N100, 
               clocked_on => CLK_port, Q => REGISTERS_53_16_port, QN => n_2711
               );
   REGISTERS_reg_53_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N125, next_state => N99, 
               clocked_on => CLK_port, Q => REGISTERS_53_15_port, QN => n_2712
               );
   REGISTERS_reg_53_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N125, next_state => N98, 
               clocked_on => CLK_port, Q => REGISTERS_53_14_port, QN => n_2713
               );
   REGISTERS_reg_53_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N125, next_state => N97, 
               clocked_on => CLK_port, Q => REGISTERS_53_13_port, QN => n_2714
               );
   REGISTERS_reg_53_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N125, next_state => N96, 
               clocked_on => CLK_port, Q => REGISTERS_53_12_port, QN => n_2715
               );
   REGISTERS_reg_53_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N125, next_state => N95, 
               clocked_on => CLK_port, Q => REGISTERS_53_11_port, QN => n_2716
               );
   REGISTERS_reg_53_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N125, next_state => N94, 
               clocked_on => CLK_port, Q => REGISTERS_53_10_port, QN => n_2717
               );
   REGISTERS_reg_53_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N125, next_state => N93, 
               clocked_on => CLK_port, Q => REGISTERS_53_9_port, QN => n_2718);
   REGISTERS_reg_53_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N125, next_state => N92, 
               clocked_on => CLK_port, Q => REGISTERS_53_8_port, QN => n_2719);
   REGISTERS_reg_53_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N125, next_state => N91, 
               clocked_on => CLK_port, Q => REGISTERS_53_7_port, QN => n_2720);
   REGISTERS_reg_53_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N125, next_state => N90, 
               clocked_on => CLK_port, Q => REGISTERS_53_6_port, QN => n_2721);
   REGISTERS_reg_53_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N125, next_state => N89, 
               clocked_on => CLK_port, Q => REGISTERS_53_5_port, QN => n_2722);
   REGISTERS_reg_53_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N125, next_state => N88, 
               clocked_on => CLK_port, Q => REGISTERS_53_4_port, QN => n_2723);
   REGISTERS_reg_53_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N125, next_state => N87, 
               clocked_on => CLK_port, Q => REGISTERS_53_3_port, QN => n_2724);
   REGISTERS_reg_53_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N125, next_state => N86, 
               clocked_on => CLK_port, Q => REGISTERS_53_2_port, QN => n_2725);
   REGISTERS_reg_53_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N125, next_state => N85, 
               clocked_on => CLK_port, Q => REGISTERS_53_1_port, QN => n_2726);
   REGISTERS_reg_53_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N125, next_state => N84, 
               clocked_on => CLK_port, Q => REGISTERS_53_0_port, QN => n_2727);
   REGISTERS_reg_54_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N124, next_state => N115, 
               clocked_on => CLK_port, Q => REGISTERS_54_31_port, QN => n_2728
               );
   REGISTERS_reg_54_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N124, next_state => N114, 
               clocked_on => CLK_port, Q => REGISTERS_54_30_port, QN => n_2729
               );
   REGISTERS_reg_54_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N124, next_state => N113, 
               clocked_on => CLK_port, Q => REGISTERS_54_29_port, QN => n_2730
               );
   REGISTERS_reg_54_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N124, next_state => N112, 
               clocked_on => CLK_port, Q => REGISTERS_54_28_port, QN => n_2731
               );
   REGISTERS_reg_54_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N124, next_state => N111, 
               clocked_on => CLK_port, Q => REGISTERS_54_27_port, QN => n_2732
               );
   REGISTERS_reg_54_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N124, next_state => N110, 
               clocked_on => CLK_port, Q => REGISTERS_54_26_port, QN => n_2733
               );
   REGISTERS_reg_54_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N124, next_state => N109, 
               clocked_on => CLK_port, Q => REGISTERS_54_25_port, QN => n_2734
               );
   REGISTERS_reg_54_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N124, next_state => N108, 
               clocked_on => CLK_port, Q => REGISTERS_54_24_port, QN => n_2735
               );
   REGISTERS_reg_54_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N124, next_state => N107, 
               clocked_on => CLK_port, Q => REGISTERS_54_23_port, QN => n_2736
               );
   REGISTERS_reg_54_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N124, next_state => N106, 
               clocked_on => CLK_port, Q => REGISTERS_54_22_port, QN => n_2737
               );
   REGISTERS_reg_54_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N124, next_state => N105, 
               clocked_on => CLK_port, Q => REGISTERS_54_21_port, QN => n_2738
               );
   REGISTERS_reg_54_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N124, next_state => N104, 
               clocked_on => CLK_port, Q => REGISTERS_54_20_port, QN => n_2739
               );
   REGISTERS_reg_54_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N124, next_state => N103, 
               clocked_on => CLK_port, Q => REGISTERS_54_19_port, QN => n_2740
               );
   REGISTERS_reg_54_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N124, next_state => N102, 
               clocked_on => CLK_port, Q => REGISTERS_54_18_port, QN => n_2741
               );
   REGISTERS_reg_54_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N124, next_state => N101, 
               clocked_on => CLK_port, Q => REGISTERS_54_17_port, QN => n_2742
               );
   REGISTERS_reg_54_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N124, next_state => N100, 
               clocked_on => CLK_port, Q => REGISTERS_54_16_port, QN => n_2743
               );
   REGISTERS_reg_54_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N124, next_state => N99, 
               clocked_on => CLK_port, Q => REGISTERS_54_15_port, QN => n_2744
               );
   REGISTERS_reg_54_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N124, next_state => N98, 
               clocked_on => CLK_port, Q => REGISTERS_54_14_port, QN => n_2745
               );
   REGISTERS_reg_54_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N124, next_state => N97, 
               clocked_on => CLK_port, Q => REGISTERS_54_13_port, QN => n_2746
               );
   REGISTERS_reg_54_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N124, next_state => N96, 
               clocked_on => CLK_port, Q => REGISTERS_54_12_port, QN => n_2747
               );
   REGISTERS_reg_54_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N124, next_state => N95, 
               clocked_on => CLK_port, Q => REGISTERS_54_11_port, QN => n_2748
               );
   REGISTERS_reg_54_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N124, next_state => N94, 
               clocked_on => CLK_port, Q => REGISTERS_54_10_port, QN => n_2749
               );
   REGISTERS_reg_54_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N124, next_state => N93, 
               clocked_on => CLK_port, Q => REGISTERS_54_9_port, QN => n_2750);
   REGISTERS_reg_54_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N124, next_state => N92, 
               clocked_on => CLK_port, Q => REGISTERS_54_8_port, QN => n_2751);
   REGISTERS_reg_54_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N124, next_state => N91, 
               clocked_on => CLK_port, Q => REGISTERS_54_7_port, QN => n_2752);
   REGISTERS_reg_54_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N124, next_state => N90, 
               clocked_on => CLK_port, Q => REGISTERS_54_6_port, QN => n_2753);
   REGISTERS_reg_54_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N124, next_state => N89, 
               clocked_on => CLK_port, Q => REGISTERS_54_5_port, QN => n_2754);
   REGISTERS_reg_54_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N124, next_state => N88, 
               clocked_on => CLK_port, Q => REGISTERS_54_4_port, QN => n_2755);
   REGISTERS_reg_54_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N124, next_state => N87, 
               clocked_on => CLK_port, Q => REGISTERS_54_3_port, QN => n_2756);
   REGISTERS_reg_54_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N124, next_state => N86, 
               clocked_on => CLK_port, Q => REGISTERS_54_2_port, QN => n_2757);
   REGISTERS_reg_54_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N124, next_state => N85, 
               clocked_on => CLK_port, Q => REGISTERS_54_1_port, QN => n_2758);
   REGISTERS_reg_54_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N124, next_state => N84, 
               clocked_on => CLK_port, Q => REGISTERS_54_0_port, QN => n_2759);
   REGISTERS_reg_55_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N123, next_state => N115, 
               clocked_on => CLK_port, Q => REGISTERS_55_31_port, QN => n_2760
               );
   REGISTERS_reg_55_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N123, next_state => N114, 
               clocked_on => CLK_port, Q => REGISTERS_55_30_port, QN => n_2761
               );
   REGISTERS_reg_55_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N123, next_state => N113, 
               clocked_on => CLK_port, Q => REGISTERS_55_29_port, QN => n_2762
               );
   REGISTERS_reg_55_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N123, next_state => N112, 
               clocked_on => CLK_port, Q => REGISTERS_55_28_port, QN => n_2763
               );
   REGISTERS_reg_55_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N123, next_state => N111, 
               clocked_on => CLK_port, Q => REGISTERS_55_27_port, QN => n_2764
               );
   REGISTERS_reg_55_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N123, next_state => N110, 
               clocked_on => CLK_port, Q => REGISTERS_55_26_port, QN => n_2765
               );
   REGISTERS_reg_55_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N123, next_state => N109, 
               clocked_on => CLK_port, Q => REGISTERS_55_25_port, QN => n_2766
               );
   REGISTERS_reg_55_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N123, next_state => N108, 
               clocked_on => CLK_port, Q => REGISTERS_55_24_port, QN => n_2767
               );
   REGISTERS_reg_55_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N123, next_state => N107, 
               clocked_on => CLK_port, Q => REGISTERS_55_23_port, QN => n_2768
               );
   REGISTERS_reg_55_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N123, next_state => N106, 
               clocked_on => CLK_port, Q => REGISTERS_55_22_port, QN => n_2769
               );
   REGISTERS_reg_55_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N123, next_state => N105, 
               clocked_on => CLK_port, Q => REGISTERS_55_21_port, QN => n_2770
               );
   REGISTERS_reg_55_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N123, next_state => N104, 
               clocked_on => CLK_port, Q => REGISTERS_55_20_port, QN => n_2771
               );
   REGISTERS_reg_55_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N123, next_state => N103, 
               clocked_on => CLK_port, Q => REGISTERS_55_19_port, QN => n_2772
               );
   REGISTERS_reg_55_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N123, next_state => N102, 
               clocked_on => CLK_port, Q => REGISTERS_55_18_port, QN => n_2773
               );
   REGISTERS_reg_55_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N123, next_state => N101, 
               clocked_on => CLK_port, Q => REGISTERS_55_17_port, QN => n_2774
               );
   REGISTERS_reg_55_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N123, next_state => N100, 
               clocked_on => CLK_port, Q => REGISTERS_55_16_port, QN => n_2775
               );
   REGISTERS_reg_55_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N123, next_state => N99, 
               clocked_on => CLK_port, Q => REGISTERS_55_15_port, QN => n_2776
               );
   REGISTERS_reg_55_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N123, next_state => N98, 
               clocked_on => CLK_port, Q => REGISTERS_55_14_port, QN => n_2777
               );
   REGISTERS_reg_55_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N123, next_state => N97, 
               clocked_on => CLK_port, Q => REGISTERS_55_13_port, QN => n_2778
               );
   REGISTERS_reg_55_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N123, next_state => N96, 
               clocked_on => CLK_port, Q => REGISTERS_55_12_port, QN => n_2779
               );
   REGISTERS_reg_55_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N123, next_state => N95, 
               clocked_on => CLK_port, Q => REGISTERS_55_11_port, QN => n_2780
               );
   REGISTERS_reg_55_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N123, next_state => N94, 
               clocked_on => CLK_port, Q => REGISTERS_55_10_port, QN => n_2781
               );
   REGISTERS_reg_55_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N123, next_state => N93, 
               clocked_on => CLK_port, Q => REGISTERS_55_9_port, QN => n_2782);
   REGISTERS_reg_55_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N123, next_state => N92, 
               clocked_on => CLK_port, Q => REGISTERS_55_8_port, QN => n_2783);
   REGISTERS_reg_55_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N123, next_state => N91, 
               clocked_on => CLK_port, Q => REGISTERS_55_7_port, QN => n_2784);
   REGISTERS_reg_55_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N123, next_state => N90, 
               clocked_on => CLK_port, Q => REGISTERS_55_6_port, QN => n_2785);
   REGISTERS_reg_55_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N123, next_state => N89, 
               clocked_on => CLK_port, Q => REGISTERS_55_5_port, QN => n_2786);
   REGISTERS_reg_55_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N123, next_state => N88, 
               clocked_on => CLK_port, Q => REGISTERS_55_4_port, QN => n_2787);
   REGISTERS_reg_55_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N123, next_state => N87, 
               clocked_on => CLK_port, Q => REGISTERS_55_3_port, QN => n_2788);
   REGISTERS_reg_55_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N123, next_state => N86, 
               clocked_on => CLK_port, Q => REGISTERS_55_2_port, QN => n_2789);
   REGISTERS_reg_55_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N123, next_state => N85, 
               clocked_on => CLK_port, Q => REGISTERS_55_1_port, QN => n_2790);
   REGISTERS_reg_55_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N123, next_state => N84, 
               clocked_on => CLK_port, Q => REGISTERS_55_0_port, QN => n_2791);
   REGISTERS_reg_56_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N122, next_state => N115, 
               clocked_on => CLK_port, Q => REGISTERS_56_31_port, QN => n_2792
               );
   REGISTERS_reg_56_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N122, next_state => N114, 
               clocked_on => CLK_port, Q => REGISTERS_56_30_port, QN => n_2793
               );
   REGISTERS_reg_56_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N122, next_state => N113, 
               clocked_on => CLK_port, Q => REGISTERS_56_29_port, QN => n_2794
               );
   REGISTERS_reg_56_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N122, next_state => N112, 
               clocked_on => CLK_port, Q => REGISTERS_56_28_port, QN => n_2795
               );
   REGISTERS_reg_56_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N122, next_state => N111, 
               clocked_on => CLK_port, Q => REGISTERS_56_27_port, QN => n_2796
               );
   REGISTERS_reg_56_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N122, next_state => N110, 
               clocked_on => CLK_port, Q => REGISTERS_56_26_port, QN => n_2797
               );
   REGISTERS_reg_56_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N122, next_state => N109, 
               clocked_on => CLK_port, Q => REGISTERS_56_25_port, QN => n_2798
               );
   REGISTERS_reg_56_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N122, next_state => N108, 
               clocked_on => CLK_port, Q => REGISTERS_56_24_port, QN => n_2799
               );
   REGISTERS_reg_56_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N122, next_state => N107, 
               clocked_on => CLK_port, Q => REGISTERS_56_23_port, QN => n_2800
               );
   REGISTERS_reg_56_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N122, next_state => N106, 
               clocked_on => CLK_port, Q => REGISTERS_56_22_port, QN => n_2801
               );
   REGISTERS_reg_56_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N122, next_state => N105, 
               clocked_on => CLK_port, Q => REGISTERS_56_21_port, QN => n_2802
               );
   REGISTERS_reg_56_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N122, next_state => N104, 
               clocked_on => CLK_port, Q => REGISTERS_56_20_port, QN => n_2803
               );
   REGISTERS_reg_56_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N122, next_state => N103, 
               clocked_on => CLK_port, Q => REGISTERS_56_19_port, QN => n_2804
               );
   REGISTERS_reg_56_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N122, next_state => N102, 
               clocked_on => CLK_port, Q => REGISTERS_56_18_port, QN => n_2805
               );
   REGISTERS_reg_56_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N122, next_state => N101, 
               clocked_on => CLK_port, Q => REGISTERS_56_17_port, QN => n_2806
               );
   REGISTERS_reg_56_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N122, next_state => N100, 
               clocked_on => CLK_port, Q => REGISTERS_56_16_port, QN => n_2807
               );
   REGISTERS_reg_56_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N122, next_state => N99, 
               clocked_on => CLK_port, Q => REGISTERS_56_15_port, QN => n_2808
               );
   REGISTERS_reg_56_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N122, next_state => N98, 
               clocked_on => CLK_port, Q => REGISTERS_56_14_port, QN => n_2809
               );
   REGISTERS_reg_56_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N122, next_state => N97, 
               clocked_on => CLK_port, Q => REGISTERS_56_13_port, QN => n_2810
               );
   REGISTERS_reg_56_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N122, next_state => N96, 
               clocked_on => CLK_port, Q => REGISTERS_56_12_port, QN => n_2811
               );
   REGISTERS_reg_56_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N122, next_state => N95, 
               clocked_on => CLK_port, Q => REGISTERS_56_11_port, QN => n_2812
               );
   REGISTERS_reg_56_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N122, next_state => N94, 
               clocked_on => CLK_port, Q => REGISTERS_56_10_port, QN => n_2813
               );
   REGISTERS_reg_56_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N122, next_state => N93, 
               clocked_on => CLK_port, Q => REGISTERS_56_9_port, QN => n_2814);
   REGISTERS_reg_56_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N122, next_state => N92, 
               clocked_on => CLK_port, Q => REGISTERS_56_8_port, QN => n_2815);
   REGISTERS_reg_56_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N122, next_state => N91, 
               clocked_on => CLK_port, Q => REGISTERS_56_7_port, QN => n_2816);
   REGISTERS_reg_56_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N122, next_state => N90, 
               clocked_on => CLK_port, Q => REGISTERS_56_6_port, QN => n_2817);
   REGISTERS_reg_56_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N122, next_state => N89, 
               clocked_on => CLK_port, Q => REGISTERS_56_5_port, QN => n_2818);
   REGISTERS_reg_56_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N122, next_state => N88, 
               clocked_on => CLK_port, Q => REGISTERS_56_4_port, QN => n_2819);
   REGISTERS_reg_56_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N122, next_state => N87, 
               clocked_on => CLK_port, Q => REGISTERS_56_3_port, QN => n_2820);
   REGISTERS_reg_56_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N122, next_state => N86, 
               clocked_on => CLK_port, Q => REGISTERS_56_2_port, QN => n_2821);
   REGISTERS_reg_56_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N122, next_state => N85, 
               clocked_on => CLK_port, Q => REGISTERS_56_1_port, QN => n_2822);
   REGISTERS_reg_56_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N122, next_state => N84, 
               clocked_on => CLK_port, Q => REGISTERS_56_0_port, QN => n_2823);
   REGISTERS_reg_57_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N121, next_state => N115, 
               clocked_on => CLK_port, Q => REGISTERS_57_31_port, QN => n_2824
               );
   REGISTERS_reg_57_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N121, next_state => N114, 
               clocked_on => CLK_port, Q => REGISTERS_57_30_port, QN => n_2825
               );
   REGISTERS_reg_57_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N121, next_state => N113, 
               clocked_on => CLK_port, Q => REGISTERS_57_29_port, QN => n_2826
               );
   REGISTERS_reg_57_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N121, next_state => N112, 
               clocked_on => CLK_port, Q => REGISTERS_57_28_port, QN => n_2827
               );
   REGISTERS_reg_57_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N121, next_state => N111, 
               clocked_on => CLK_port, Q => REGISTERS_57_27_port, QN => n_2828
               );
   REGISTERS_reg_57_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N121, next_state => N110, 
               clocked_on => CLK_port, Q => REGISTERS_57_26_port, QN => n_2829
               );
   REGISTERS_reg_57_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N121, next_state => N109, 
               clocked_on => CLK_port, Q => REGISTERS_57_25_port, QN => n_2830
               );
   REGISTERS_reg_57_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N121, next_state => N108, 
               clocked_on => CLK_port, Q => REGISTERS_57_24_port, QN => n_2831
               );
   REGISTERS_reg_57_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N121, next_state => N107, 
               clocked_on => CLK_port, Q => REGISTERS_57_23_port, QN => n_2832
               );
   REGISTERS_reg_57_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N121, next_state => N106, 
               clocked_on => CLK_port, Q => REGISTERS_57_22_port, QN => n_2833
               );
   REGISTERS_reg_57_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N121, next_state => N105, 
               clocked_on => CLK_port, Q => REGISTERS_57_21_port, QN => n_2834
               );
   REGISTERS_reg_57_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N121, next_state => N104, 
               clocked_on => CLK_port, Q => REGISTERS_57_20_port, QN => n_2835
               );
   REGISTERS_reg_57_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N121, next_state => N103, 
               clocked_on => CLK_port, Q => REGISTERS_57_19_port, QN => n_2836
               );
   REGISTERS_reg_57_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N121, next_state => N102, 
               clocked_on => CLK_port, Q => REGISTERS_57_18_port, QN => n_2837
               );
   REGISTERS_reg_57_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N121, next_state => N101, 
               clocked_on => CLK_port, Q => REGISTERS_57_17_port, QN => n_2838
               );
   REGISTERS_reg_57_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N121, next_state => N100, 
               clocked_on => CLK_port, Q => REGISTERS_57_16_port, QN => n_2839
               );
   REGISTERS_reg_57_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N121, next_state => N99, 
               clocked_on => CLK_port, Q => REGISTERS_57_15_port, QN => n_2840
               );
   REGISTERS_reg_57_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N121, next_state => N98, 
               clocked_on => CLK_port, Q => REGISTERS_57_14_port, QN => n_2841
               );
   REGISTERS_reg_57_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N121, next_state => N97, 
               clocked_on => CLK_port, Q => REGISTERS_57_13_port, QN => n_2842
               );
   REGISTERS_reg_57_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N121, next_state => N96, 
               clocked_on => CLK_port, Q => REGISTERS_57_12_port, QN => n_2843
               );
   REGISTERS_reg_57_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N121, next_state => N95, 
               clocked_on => CLK_port, Q => REGISTERS_57_11_port, QN => n_2844
               );
   REGISTERS_reg_57_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N121, next_state => N94, 
               clocked_on => CLK_port, Q => REGISTERS_57_10_port, QN => n_2845
               );
   REGISTERS_reg_57_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N121, next_state => N93, 
               clocked_on => CLK_port, Q => REGISTERS_57_9_port, QN => n_2846);
   REGISTERS_reg_57_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N121, next_state => N92, 
               clocked_on => CLK_port, Q => REGISTERS_57_8_port, QN => n_2847);
   REGISTERS_reg_57_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N121, next_state => N91, 
               clocked_on => CLK_port, Q => REGISTERS_57_7_port, QN => n_2848);
   REGISTERS_reg_57_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N121, next_state => N90, 
               clocked_on => CLK_port, Q => REGISTERS_57_6_port, QN => n_2849);
   REGISTERS_reg_57_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N121, next_state => N89, 
               clocked_on => CLK_port, Q => REGISTERS_57_5_port, QN => n_2850);
   REGISTERS_reg_57_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N121, next_state => N88, 
               clocked_on => CLK_port, Q => REGISTERS_57_4_port, QN => n_2851);
   REGISTERS_reg_57_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N121, next_state => N87, 
               clocked_on => CLK_port, Q => REGISTERS_57_3_port, QN => n_2852);
   REGISTERS_reg_57_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N121, next_state => N86, 
               clocked_on => CLK_port, Q => REGISTERS_57_2_port, QN => n_2853);
   REGISTERS_reg_57_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N121, next_state => N85, 
               clocked_on => CLK_port, Q => REGISTERS_57_1_port, QN => n_2854);
   REGISTERS_reg_57_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N121, next_state => N84, 
               clocked_on => CLK_port, Q => REGISTERS_57_0_port, QN => n_2855);
   REGISTERS_reg_58_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N120, next_state => N115, 
               clocked_on => CLK_port, Q => REGISTERS_58_31_port, QN => n_2856
               );
   REGISTERS_reg_58_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N120, next_state => N114, 
               clocked_on => CLK_port, Q => REGISTERS_58_30_port, QN => n_2857
               );
   REGISTERS_reg_58_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N120, next_state => N113, 
               clocked_on => CLK_port, Q => REGISTERS_58_29_port, QN => n_2858
               );
   REGISTERS_reg_58_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N120, next_state => N112, 
               clocked_on => CLK_port, Q => REGISTERS_58_28_port, QN => n_2859
               );
   REGISTERS_reg_58_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N120, next_state => N111, 
               clocked_on => CLK_port, Q => REGISTERS_58_27_port, QN => n_2860
               );
   REGISTERS_reg_58_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N120, next_state => N110, 
               clocked_on => CLK_port, Q => REGISTERS_58_26_port, QN => n_2861
               );
   REGISTERS_reg_58_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N120, next_state => N109, 
               clocked_on => CLK_port, Q => REGISTERS_58_25_port, QN => n_2862
               );
   REGISTERS_reg_58_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N120, next_state => N108, 
               clocked_on => CLK_port, Q => REGISTERS_58_24_port, QN => n_2863
               );
   REGISTERS_reg_58_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N120, next_state => N107, 
               clocked_on => CLK_port, Q => REGISTERS_58_23_port, QN => n_2864
               );
   REGISTERS_reg_58_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N120, next_state => N106, 
               clocked_on => CLK_port, Q => REGISTERS_58_22_port, QN => n_2865
               );
   REGISTERS_reg_58_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N120, next_state => N105, 
               clocked_on => CLK_port, Q => REGISTERS_58_21_port, QN => n_2866
               );
   REGISTERS_reg_58_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N120, next_state => N104, 
               clocked_on => CLK_port, Q => REGISTERS_58_20_port, QN => n_2867
               );
   REGISTERS_reg_58_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N120, next_state => N103, 
               clocked_on => CLK_port, Q => REGISTERS_58_19_port, QN => n_2868
               );
   REGISTERS_reg_58_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N120, next_state => N102, 
               clocked_on => CLK_port, Q => REGISTERS_58_18_port, QN => n_2869
               );
   REGISTERS_reg_58_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N120, next_state => N101, 
               clocked_on => CLK_port, Q => REGISTERS_58_17_port, QN => n_2870
               );
   REGISTERS_reg_58_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N120, next_state => N100, 
               clocked_on => CLK_port, Q => REGISTERS_58_16_port, QN => n_2871
               );
   REGISTERS_reg_58_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N120, next_state => N99, 
               clocked_on => CLK_port, Q => REGISTERS_58_15_port, QN => n_2872
               );
   REGISTERS_reg_58_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N120, next_state => N98, 
               clocked_on => CLK_port, Q => REGISTERS_58_14_port, QN => n_2873
               );
   REGISTERS_reg_58_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N120, next_state => N97, 
               clocked_on => CLK_port, Q => REGISTERS_58_13_port, QN => n_2874
               );
   REGISTERS_reg_58_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N120, next_state => N96, 
               clocked_on => CLK_port, Q => REGISTERS_58_12_port, QN => n_2875
               );
   REGISTERS_reg_58_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N120, next_state => N95, 
               clocked_on => CLK_port, Q => REGISTERS_58_11_port, QN => n_2876
               );
   REGISTERS_reg_58_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N120, next_state => N94, 
               clocked_on => CLK_port, Q => REGISTERS_58_10_port, QN => n_2877
               );
   REGISTERS_reg_58_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N120, next_state => N93, 
               clocked_on => CLK_port, Q => REGISTERS_58_9_port, QN => n_2878);
   REGISTERS_reg_58_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N120, next_state => N92, 
               clocked_on => CLK_port, Q => REGISTERS_58_8_port, QN => n_2879);
   REGISTERS_reg_58_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N120, next_state => N91, 
               clocked_on => CLK_port, Q => REGISTERS_58_7_port, QN => n_2880);
   REGISTERS_reg_58_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N120, next_state => N90, 
               clocked_on => CLK_port, Q => REGISTERS_58_6_port, QN => n_2881);
   REGISTERS_reg_58_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N120, next_state => N89, 
               clocked_on => CLK_port, Q => REGISTERS_58_5_port, QN => n_2882);
   REGISTERS_reg_58_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N120, next_state => N88, 
               clocked_on => CLK_port, Q => REGISTERS_58_4_port, QN => n_2883);
   REGISTERS_reg_58_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N120, next_state => N87, 
               clocked_on => CLK_port, Q => REGISTERS_58_3_port, QN => n_2884);
   REGISTERS_reg_58_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N120, next_state => N86, 
               clocked_on => CLK_port, Q => REGISTERS_58_2_port, QN => n_2885);
   REGISTERS_reg_58_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N120, next_state => N85, 
               clocked_on => CLK_port, Q => REGISTERS_58_1_port, QN => n_2886);
   REGISTERS_reg_58_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N120, next_state => N84, 
               clocked_on => CLK_port, Q => REGISTERS_58_0_port, QN => n_2887);
   REGISTERS_reg_59_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N119, next_state => N115, 
               clocked_on => CLK_port, Q => REGISTERS_59_31_port, QN => n_2888
               );
   REGISTERS_reg_59_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N119, next_state => N114, 
               clocked_on => CLK_port, Q => REGISTERS_59_30_port, QN => n_2889
               );
   REGISTERS_reg_59_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N119, next_state => N113, 
               clocked_on => CLK_port, Q => REGISTERS_59_29_port, QN => n_2890
               );
   REGISTERS_reg_59_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N119, next_state => N112, 
               clocked_on => CLK_port, Q => REGISTERS_59_28_port, QN => n_2891
               );
   REGISTERS_reg_59_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N119, next_state => N111, 
               clocked_on => CLK_port, Q => REGISTERS_59_27_port, QN => n_2892
               );
   REGISTERS_reg_59_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N119, next_state => N110, 
               clocked_on => CLK_port, Q => REGISTERS_59_26_port, QN => n_2893
               );
   REGISTERS_reg_59_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N119, next_state => N109, 
               clocked_on => CLK_port, Q => REGISTERS_59_25_port, QN => n_2894
               );
   REGISTERS_reg_59_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N119, next_state => N108, 
               clocked_on => CLK_port, Q => REGISTERS_59_24_port, QN => n_2895
               );
   REGISTERS_reg_59_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N119, next_state => N107, 
               clocked_on => CLK_port, Q => REGISTERS_59_23_port, QN => n_2896
               );
   REGISTERS_reg_59_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N119, next_state => N106, 
               clocked_on => CLK_port, Q => REGISTERS_59_22_port, QN => n_2897
               );
   REGISTERS_reg_59_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N119, next_state => N105, 
               clocked_on => CLK_port, Q => REGISTERS_59_21_port, QN => n_2898
               );
   REGISTERS_reg_59_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N119, next_state => N104, 
               clocked_on => CLK_port, Q => REGISTERS_59_20_port, QN => n_2899
               );
   REGISTERS_reg_59_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N119, next_state => N103, 
               clocked_on => CLK_port, Q => REGISTERS_59_19_port, QN => n_2900
               );
   REGISTERS_reg_59_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N119, next_state => N102, 
               clocked_on => CLK_port, Q => REGISTERS_59_18_port, QN => n_2901
               );
   REGISTERS_reg_59_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N119, next_state => N101, 
               clocked_on => CLK_port, Q => REGISTERS_59_17_port, QN => n_2902
               );
   REGISTERS_reg_59_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N119, next_state => N100, 
               clocked_on => CLK_port, Q => REGISTERS_59_16_port, QN => n_2903
               );
   REGISTERS_reg_59_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N119, next_state => N99, 
               clocked_on => CLK_port, Q => REGISTERS_59_15_port, QN => n_2904
               );
   REGISTERS_reg_59_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N119, next_state => N98, 
               clocked_on => CLK_port, Q => REGISTERS_59_14_port, QN => n_2905
               );
   REGISTERS_reg_59_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N119, next_state => N97, 
               clocked_on => CLK_port, Q => REGISTERS_59_13_port, QN => n_2906
               );
   REGISTERS_reg_59_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N119, next_state => N96, 
               clocked_on => CLK_port, Q => REGISTERS_59_12_port, QN => n_2907
               );
   REGISTERS_reg_59_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N119, next_state => N95, 
               clocked_on => CLK_port, Q => REGISTERS_59_11_port, QN => n_2908
               );
   REGISTERS_reg_59_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N119, next_state => N94, 
               clocked_on => CLK_port, Q => REGISTERS_59_10_port, QN => n_2909
               );
   REGISTERS_reg_59_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N119, next_state => N93, 
               clocked_on => CLK_port, Q => REGISTERS_59_9_port, QN => n_2910);
   REGISTERS_reg_59_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N119, next_state => N92, 
               clocked_on => CLK_port, Q => REGISTERS_59_8_port, QN => n_2911);
   REGISTERS_reg_59_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N119, next_state => N91, 
               clocked_on => CLK_port, Q => REGISTERS_59_7_port, QN => n_2912);
   REGISTERS_reg_59_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N119, next_state => N90, 
               clocked_on => CLK_port, Q => REGISTERS_59_6_port, QN => n_2913);
   REGISTERS_reg_59_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N119, next_state => N89, 
               clocked_on => CLK_port, Q => REGISTERS_59_5_port, QN => n_2914);
   REGISTERS_reg_59_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N119, next_state => N88, 
               clocked_on => CLK_port, Q => REGISTERS_59_4_port, QN => n_2915);
   REGISTERS_reg_59_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N119, next_state => N87, 
               clocked_on => CLK_port, Q => REGISTERS_59_3_port, QN => n_2916);
   REGISTERS_reg_59_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N119, next_state => N86, 
               clocked_on => CLK_port, Q => REGISTERS_59_2_port, QN => n_2917);
   REGISTERS_reg_59_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N119, next_state => N85, 
               clocked_on => CLK_port, Q => REGISTERS_59_1_port, QN => n_2918);
   REGISTERS_reg_59_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N119, next_state => N84, 
               clocked_on => CLK_port, Q => REGISTERS_59_0_port, QN => n_2919);
   REGISTERS_reg_60_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N118, next_state => N115, 
               clocked_on => CLK_port, Q => REGISTERS_60_31_port, QN => n_2920
               );
   REGISTERS_reg_60_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N118, next_state => N114, 
               clocked_on => CLK_port, Q => REGISTERS_60_30_port, QN => n_2921
               );
   REGISTERS_reg_60_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N118, next_state => N113, 
               clocked_on => CLK_port, Q => REGISTERS_60_29_port, QN => n_2922
               );
   REGISTERS_reg_60_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N118, next_state => N112, 
               clocked_on => CLK_port, Q => REGISTERS_60_28_port, QN => n_2923
               );
   REGISTERS_reg_60_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N118, next_state => N111, 
               clocked_on => CLK_port, Q => REGISTERS_60_27_port, QN => n_2924
               );
   REGISTERS_reg_60_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N118, next_state => N110, 
               clocked_on => CLK_port, Q => REGISTERS_60_26_port, QN => n_2925
               );
   REGISTERS_reg_60_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N118, next_state => N109, 
               clocked_on => CLK_port, Q => REGISTERS_60_25_port, QN => n_2926
               );
   REGISTERS_reg_60_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N118, next_state => N108, 
               clocked_on => CLK_port, Q => REGISTERS_60_24_port, QN => n_2927
               );
   REGISTERS_reg_60_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N118, next_state => N107, 
               clocked_on => CLK_port, Q => REGISTERS_60_23_port, QN => n_2928
               );
   REGISTERS_reg_60_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N118, next_state => N106, 
               clocked_on => CLK_port, Q => REGISTERS_60_22_port, QN => n_2929
               );
   REGISTERS_reg_60_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N118, next_state => N105, 
               clocked_on => CLK_port, Q => REGISTERS_60_21_port, QN => n_2930
               );
   REGISTERS_reg_60_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N118, next_state => N104, 
               clocked_on => CLK_port, Q => REGISTERS_60_20_port, QN => n_2931
               );
   REGISTERS_reg_60_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N118, next_state => N103, 
               clocked_on => CLK_port, Q => REGISTERS_60_19_port, QN => n_2932
               );
   REGISTERS_reg_60_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N118, next_state => N102, 
               clocked_on => CLK_port, Q => REGISTERS_60_18_port, QN => n_2933
               );
   REGISTERS_reg_60_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N118, next_state => N101, 
               clocked_on => CLK_port, Q => REGISTERS_60_17_port, QN => n_2934
               );
   REGISTERS_reg_60_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N118, next_state => N100, 
               clocked_on => CLK_port, Q => REGISTERS_60_16_port, QN => n_2935
               );
   REGISTERS_reg_60_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N118, next_state => N99, 
               clocked_on => CLK_port, Q => REGISTERS_60_15_port, QN => n_2936
               );
   REGISTERS_reg_60_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N118, next_state => N98, 
               clocked_on => CLK_port, Q => REGISTERS_60_14_port, QN => n_2937
               );
   REGISTERS_reg_60_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N118, next_state => N97, 
               clocked_on => CLK_port, Q => REGISTERS_60_13_port, QN => n_2938
               );
   REGISTERS_reg_60_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N118, next_state => N96, 
               clocked_on => CLK_port, Q => REGISTERS_60_12_port, QN => n_2939
               );
   REGISTERS_reg_60_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N118, next_state => N95, 
               clocked_on => CLK_port, Q => REGISTERS_60_11_port, QN => n_2940
               );
   REGISTERS_reg_60_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N118, next_state => N94, 
               clocked_on => CLK_port, Q => REGISTERS_60_10_port, QN => n_2941
               );
   REGISTERS_reg_60_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N118, next_state => N93, 
               clocked_on => CLK_port, Q => REGISTERS_60_9_port, QN => n_2942);
   REGISTERS_reg_60_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N118, next_state => N92, 
               clocked_on => CLK_port, Q => REGISTERS_60_8_port, QN => n_2943);
   REGISTERS_reg_60_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N118, next_state => N91, 
               clocked_on => CLK_port, Q => REGISTERS_60_7_port, QN => n_2944);
   REGISTERS_reg_60_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N118, next_state => N90, 
               clocked_on => CLK_port, Q => REGISTERS_60_6_port, QN => n_2945);
   REGISTERS_reg_60_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N118, next_state => N89, 
               clocked_on => CLK_port, Q => REGISTERS_60_5_port, QN => n_2946);
   REGISTERS_reg_60_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N118, next_state => N88, 
               clocked_on => CLK_port, Q => REGISTERS_60_4_port, QN => n_2947);
   REGISTERS_reg_60_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N118, next_state => N87, 
               clocked_on => CLK_port, Q => REGISTERS_60_3_port, QN => n_2948);
   REGISTERS_reg_60_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N118, next_state => N86, 
               clocked_on => CLK_port, Q => REGISTERS_60_2_port, QN => n_2949);
   REGISTERS_reg_60_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N118, next_state => N85, 
               clocked_on => CLK_port, Q => REGISTERS_60_1_port, QN => n_2950);
   REGISTERS_reg_60_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N118, next_state => N84, 
               clocked_on => CLK_port, Q => REGISTERS_60_0_port, QN => n_2951);
   REGISTERS_reg_61_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N117, next_state => N115, 
               clocked_on => CLK_port, Q => REGISTERS_61_31_port, QN => n_2952
               );
   REGISTERS_reg_61_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N117, next_state => N114, 
               clocked_on => CLK_port, Q => REGISTERS_61_30_port, QN => n_2953
               );
   REGISTERS_reg_61_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N117, next_state => N113, 
               clocked_on => CLK_port, Q => REGISTERS_61_29_port, QN => n_2954
               );
   REGISTERS_reg_61_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N117, next_state => N112, 
               clocked_on => CLK_port, Q => REGISTERS_61_28_port, QN => n_2955
               );
   REGISTERS_reg_61_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N117, next_state => N111, 
               clocked_on => CLK_port, Q => REGISTERS_61_27_port, QN => n_2956
               );
   REGISTERS_reg_61_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N117, next_state => N110, 
               clocked_on => CLK_port, Q => REGISTERS_61_26_port, QN => n_2957
               );
   REGISTERS_reg_61_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N117, next_state => N109, 
               clocked_on => CLK_port, Q => REGISTERS_61_25_port, QN => n_2958
               );
   REGISTERS_reg_61_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N117, next_state => N108, 
               clocked_on => CLK_port, Q => REGISTERS_61_24_port, QN => n_2959
               );
   REGISTERS_reg_61_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N117, next_state => N107, 
               clocked_on => CLK_port, Q => REGISTERS_61_23_port, QN => n_2960
               );
   REGISTERS_reg_61_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N117, next_state => N106, 
               clocked_on => CLK_port, Q => REGISTERS_61_22_port, QN => n_2961
               );
   REGISTERS_reg_61_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N117, next_state => N105, 
               clocked_on => CLK_port, Q => REGISTERS_61_21_port, QN => n_2962
               );
   REGISTERS_reg_61_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N117, next_state => N104, 
               clocked_on => CLK_port, Q => REGISTERS_61_20_port, QN => n_2963
               );
   REGISTERS_reg_61_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N117, next_state => N103, 
               clocked_on => CLK_port, Q => REGISTERS_61_19_port, QN => n_2964
               );
   REGISTERS_reg_61_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N117, next_state => N102, 
               clocked_on => CLK_port, Q => REGISTERS_61_18_port, QN => n_2965
               );
   REGISTERS_reg_61_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N117, next_state => N101, 
               clocked_on => CLK_port, Q => REGISTERS_61_17_port, QN => n_2966
               );
   REGISTERS_reg_61_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N117, next_state => N100, 
               clocked_on => CLK_port, Q => REGISTERS_61_16_port, QN => n_2967
               );
   REGISTERS_reg_61_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N117, next_state => N99, 
               clocked_on => CLK_port, Q => REGISTERS_61_15_port, QN => n_2968
               );
   REGISTERS_reg_61_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N117, next_state => N98, 
               clocked_on => CLK_port, Q => REGISTERS_61_14_port, QN => n_2969
               );
   REGISTERS_reg_61_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N117, next_state => N97, 
               clocked_on => CLK_port, Q => REGISTERS_61_13_port, QN => n_2970
               );
   REGISTERS_reg_61_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N117, next_state => N96, 
               clocked_on => CLK_port, Q => REGISTERS_61_12_port, QN => n_2971
               );
   REGISTERS_reg_61_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N117, next_state => N95, 
               clocked_on => CLK_port, Q => REGISTERS_61_11_port, QN => n_2972
               );
   REGISTERS_reg_61_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N117, next_state => N94, 
               clocked_on => CLK_port, Q => REGISTERS_61_10_port, QN => n_2973
               );
   REGISTERS_reg_61_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N117, next_state => N93, 
               clocked_on => CLK_port, Q => REGISTERS_61_9_port, QN => n_2974);
   REGISTERS_reg_61_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N117, next_state => N92, 
               clocked_on => CLK_port, Q => REGISTERS_61_8_port, QN => n_2975);
   REGISTERS_reg_61_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N117, next_state => N91, 
               clocked_on => CLK_port, Q => REGISTERS_61_7_port, QN => n_2976);
   REGISTERS_reg_61_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N117, next_state => N90, 
               clocked_on => CLK_port, Q => REGISTERS_61_6_port, QN => n_2977);
   REGISTERS_reg_61_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N117, next_state => N89, 
               clocked_on => CLK_port, Q => REGISTERS_61_5_port, QN => n_2978);
   REGISTERS_reg_61_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N117, next_state => N88, 
               clocked_on => CLK_port, Q => REGISTERS_61_4_port, QN => n_2979);
   REGISTERS_reg_61_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N117, next_state => N87, 
               clocked_on => CLK_port, Q => REGISTERS_61_3_port, QN => n_2980);
   REGISTERS_reg_61_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N117, next_state => N86, 
               clocked_on => CLK_port, Q => REGISTERS_61_2_port, QN => n_2981);
   REGISTERS_reg_61_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N117, next_state => N85, 
               clocked_on => CLK_port, Q => REGISTERS_61_1_port, QN => n_2982);
   REGISTERS_reg_61_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N117, next_state => N84, 
               clocked_on => CLK_port, Q => REGISTERS_61_0_port, QN => n_2983);
   REGISTERS_reg_62_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N116, next_state => N115, 
               clocked_on => CLK_port, Q => REGISTERS_62_31_port, QN => n_2984
               );
   REGISTERS_reg_62_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N116, next_state => N114, 
               clocked_on => CLK_port, Q => REGISTERS_62_30_port, QN => n_2985
               );
   REGISTERS_reg_62_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N116, next_state => N113, 
               clocked_on => CLK_port, Q => REGISTERS_62_29_port, QN => n_2986
               );
   REGISTERS_reg_62_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N116, next_state => N112, 
               clocked_on => CLK_port, Q => REGISTERS_62_28_port, QN => n_2987
               );
   REGISTERS_reg_62_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N116, next_state => N111, 
               clocked_on => CLK_port, Q => REGISTERS_62_27_port, QN => n_2988
               );
   REGISTERS_reg_62_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N116, next_state => N110, 
               clocked_on => CLK_port, Q => REGISTERS_62_26_port, QN => n_2989
               );
   REGISTERS_reg_62_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N116, next_state => N109, 
               clocked_on => CLK_port, Q => REGISTERS_62_25_port, QN => n_2990
               );
   REGISTERS_reg_62_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N116, next_state => N108, 
               clocked_on => CLK_port, Q => REGISTERS_62_24_port, QN => n_2991
               );
   REGISTERS_reg_62_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N116, next_state => N107, 
               clocked_on => CLK_port, Q => REGISTERS_62_23_port, QN => n_2992
               );
   REGISTERS_reg_62_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N116, next_state => N106, 
               clocked_on => CLK_port, Q => REGISTERS_62_22_port, QN => n_2993
               );
   REGISTERS_reg_62_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N116, next_state => N105, 
               clocked_on => CLK_port, Q => REGISTERS_62_21_port, QN => n_2994
               );
   REGISTERS_reg_62_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N116, next_state => N104, 
               clocked_on => CLK_port, Q => REGISTERS_62_20_port, QN => n_2995
               );
   REGISTERS_reg_62_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N116, next_state => N103, 
               clocked_on => CLK_port, Q => REGISTERS_62_19_port, QN => n_2996
               );
   REGISTERS_reg_62_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N116, next_state => N102, 
               clocked_on => CLK_port, Q => REGISTERS_62_18_port, QN => n_2997
               );
   REGISTERS_reg_62_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N116, next_state => N101, 
               clocked_on => CLK_port, Q => REGISTERS_62_17_port, QN => n_2998
               );
   REGISTERS_reg_62_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N116, next_state => N100, 
               clocked_on => CLK_port, Q => REGISTERS_62_16_port, QN => n_2999
               );
   REGISTERS_reg_62_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N116, next_state => N99, 
               clocked_on => CLK_port, Q => REGISTERS_62_15_port, QN => n_3000
               );
   REGISTERS_reg_62_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N116, next_state => N98, 
               clocked_on => CLK_port, Q => REGISTERS_62_14_port, QN => n_3001
               );
   REGISTERS_reg_62_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N116, next_state => N97, 
               clocked_on => CLK_port, Q => REGISTERS_62_13_port, QN => n_3002
               );
   REGISTERS_reg_62_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N116, next_state => N96, 
               clocked_on => CLK_port, Q => REGISTERS_62_12_port, QN => n_3003
               );
   REGISTERS_reg_62_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N116, next_state => N95, 
               clocked_on => CLK_port, Q => REGISTERS_62_11_port, QN => n_3004
               );
   REGISTERS_reg_62_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N116, next_state => N94, 
               clocked_on => CLK_port, Q => REGISTERS_62_10_port, QN => n_3005
               );
   REGISTERS_reg_62_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N116, next_state => N93, 
               clocked_on => CLK_port, Q => REGISTERS_62_9_port, QN => n_3006);
   REGISTERS_reg_62_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N116, next_state => N92, 
               clocked_on => CLK_port, Q => REGISTERS_62_8_port, QN => n_3007);
   REGISTERS_reg_62_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N116, next_state => N91, 
               clocked_on => CLK_port, Q => REGISTERS_62_7_port, QN => n_3008);
   REGISTERS_reg_62_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N116, next_state => N90, 
               clocked_on => CLK_port, Q => REGISTERS_62_6_port, QN => n_3009);
   REGISTERS_reg_62_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N116, next_state => N89, 
               clocked_on => CLK_port, Q => REGISTERS_62_5_port, QN => n_3010);
   REGISTERS_reg_62_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N116, next_state => N88, 
               clocked_on => CLK_port, Q => REGISTERS_62_4_port, QN => n_3011);
   REGISTERS_reg_62_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N116, next_state => N87, 
               clocked_on => CLK_port, Q => REGISTERS_62_3_port, QN => n_3012);
   REGISTERS_reg_62_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N116, next_state => N86, 
               clocked_on => CLK_port, Q => REGISTERS_62_2_port, QN => n_3013);
   REGISTERS_reg_62_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N116, next_state => N85, 
               clocked_on => CLK_port, Q => REGISTERS_62_1_port, QN => n_3014);
   REGISTERS_reg_62_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N116, next_state => N84, 
               clocked_on => CLK_port, Q => REGISTERS_62_0_port, QN => n_3015);
   REGISTERS_reg_63_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N83, next_state => N115, 
               clocked_on => CLK_port, Q => REGISTERS_63_31_port, QN => n_3016
               );
   REGISTERS_reg_63_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N83, next_state => N114, 
               clocked_on => CLK_port, Q => REGISTERS_63_30_port, QN => n_3017
               );
   REGISTERS_reg_63_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N83, next_state => N113, 
               clocked_on => CLK_port, Q => REGISTERS_63_29_port, QN => n_3018
               );
   REGISTERS_reg_63_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N83, next_state => N112, 
               clocked_on => CLK_port, Q => REGISTERS_63_28_port, QN => n_3019
               );
   REGISTERS_reg_63_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N83, next_state => N111, 
               clocked_on => CLK_port, Q => REGISTERS_63_27_port, QN => n_3020
               );
   REGISTERS_reg_63_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N83, next_state => N110, 
               clocked_on => CLK_port, Q => REGISTERS_63_26_port, QN => n_3021
               );
   REGISTERS_reg_63_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N83, next_state => N109, 
               clocked_on => CLK_port, Q => REGISTERS_63_25_port, QN => n_3022
               );
   REGISTERS_reg_63_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N83, next_state => N108, 
               clocked_on => CLK_port, Q => REGISTERS_63_24_port, QN => n_3023
               );
   REGISTERS_reg_63_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N83, next_state => N107, 
               clocked_on => CLK_port, Q => REGISTERS_63_23_port, QN => n_3024
               );
   REGISTERS_reg_63_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N83, next_state => N106, 
               clocked_on => CLK_port, Q => REGISTERS_63_22_port, QN => n_3025
               );
   REGISTERS_reg_63_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N83, next_state => N105, 
               clocked_on => CLK_port, Q => REGISTERS_63_21_port, QN => n_3026
               );
   REGISTERS_reg_63_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N83, next_state => N104, 
               clocked_on => CLK_port, Q => REGISTERS_63_20_port, QN => n_3027
               );
   REGISTERS_reg_63_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N83, next_state => N103, 
               clocked_on => CLK_port, Q => REGISTERS_63_19_port, QN => n_3028
               );
   REGISTERS_reg_63_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N83, next_state => N102, 
               clocked_on => CLK_port, Q => REGISTERS_63_18_port, QN => n_3029
               );
   REGISTERS_reg_63_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N83, next_state => N101, 
               clocked_on => CLK_port, Q => REGISTERS_63_17_port, QN => n_3030
               );
   REGISTERS_reg_63_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N83, next_state => N100, 
               clocked_on => CLK_port, Q => REGISTERS_63_16_port, QN => n_3031
               );
   REGISTERS_reg_63_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N83, next_state => N99, 
               clocked_on => CLK_port, Q => REGISTERS_63_15_port, QN => n_3032
               );
   REGISTERS_reg_63_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N83, next_state => N98, 
               clocked_on => CLK_port, Q => REGISTERS_63_14_port, QN => n_3033
               );
   REGISTERS_reg_63_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N83, next_state => N97, 
               clocked_on => CLK_port, Q => REGISTERS_63_13_port, QN => n_3034
               );
   REGISTERS_reg_63_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N83, next_state => N96, 
               clocked_on => CLK_port, Q => REGISTERS_63_12_port, QN => n_3035
               );
   REGISTERS_reg_63_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N83, next_state => N95, 
               clocked_on => CLK_port, Q => REGISTERS_63_11_port, QN => n_3036
               );
   REGISTERS_reg_63_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N83, next_state => N94, 
               clocked_on => CLK_port, Q => REGISTERS_63_10_port, QN => n_3037
               );
   REGISTERS_reg_63_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N83, next_state => N93, 
               clocked_on => CLK_port, Q => REGISTERS_63_9_port, QN => n_3038);
   REGISTERS_reg_63_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N83, next_state => N92, 
               clocked_on => CLK_port, Q => REGISTERS_63_8_port, QN => n_3039);
   REGISTERS_reg_63_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N83, next_state => N91, 
               clocked_on => CLK_port, Q => REGISTERS_63_7_port, QN => n_3040);
   REGISTERS_reg_63_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N83, next_state => N90, 
               clocked_on => CLK_port, Q => REGISTERS_63_6_port, QN => n_3041);
   REGISTERS_reg_63_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N83, next_state => N89, 
               clocked_on => CLK_port, Q => REGISTERS_63_5_port, QN => n_3042);
   REGISTERS_reg_63_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N83, next_state => N88, 
               clocked_on => CLK_port, Q => REGISTERS_63_4_port, QN => n_3043);
   REGISTERS_reg_63_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N83, next_state => N87, 
               clocked_on => CLK_port, Q => REGISTERS_63_3_port, QN => n_3044);
   REGISTERS_reg_63_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N83, next_state => N86, 
               clocked_on => CLK_port, Q => REGISTERS_63_2_port, QN => n_3045);
   REGISTERS_reg_63_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N83, next_state => N85, 
               clocked_on => CLK_port, Q => REGISTERS_63_1_port, QN => n_3046);
   REGISTERS_reg_63_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N83, next_state => N84, 
               clocked_on => CLK_port, Q => REGISTERS_63_0_port, QN => n_3047);
   C12729_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_31_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_31_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_31_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_31_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_31_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_31_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_31_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_31_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_31_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_31_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_31_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_31_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_31_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_31_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_31_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_31_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_31_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_31_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_31_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_31_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_31_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_31_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_31_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_31_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_31_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_31_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_31_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_31_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_31_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_31_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_31_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_31_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_31_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_31_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_31_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_31_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_31_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_31_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_31_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_31_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_31_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_31_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_31_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_31_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_31_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_31_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_31_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_31_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_31_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_31_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_31_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_31_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_31_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_31_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_31_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_31_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_31_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_31_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_31_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_31_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_31_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_31_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_31_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_31_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N248, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N252, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N254, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N256, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N258, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N260, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N262, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N264, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N266, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N268, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N270, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N272, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N274, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N276, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N278, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N280, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N282, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N284, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N286, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N288, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N290, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N292, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N294, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N296, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N298, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N300, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N302, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N304, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N306, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N308, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N310, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N249, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N251, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N253, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N255, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N257, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N259, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N261, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N263, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N265, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N267, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N269, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N271, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N273, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N275, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N277, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N279, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N281, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N283, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N285, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N287, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N289, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N291, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N293, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N295, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N297, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N299, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N301, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N303, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N305, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N307, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N309, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N311, 
         -- Connections to port 'Z'
         Z(0) => N312 );
   C12730_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_30_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_30_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_30_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_30_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_30_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_30_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_30_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_30_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_30_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_30_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_30_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_30_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_30_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_30_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_30_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_30_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_30_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_30_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_30_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_30_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_30_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_30_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_30_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_30_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_30_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_30_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_30_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_30_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_30_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_30_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_30_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_30_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_30_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_30_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_30_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_30_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_30_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_30_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_30_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_30_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_30_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_30_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_30_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_30_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_30_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_30_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_30_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_30_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_30_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_30_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_30_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_30_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_30_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_30_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_30_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_30_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_30_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_30_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_30_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_30_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_30_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_30_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_30_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_30_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N248, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N252, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N254, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N256, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N258, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N260, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N262, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N264, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N266, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N268, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N270, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N272, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N274, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N276, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N278, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N280, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N282, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N284, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N286, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N288, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N290, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N292, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N294, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N296, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N298, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N300, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N302, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N304, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N306, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N308, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N310, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N249, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N251, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N253, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N255, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N257, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N259, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N261, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N263, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N265, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N267, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N269, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N271, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N273, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N275, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N277, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N279, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N281, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N283, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N285, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N287, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N289, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N291, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N293, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N295, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N297, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N299, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N301, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N303, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N305, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N307, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N309, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N311, 
         -- Connections to port 'Z'
         Z(0) => N313 );
   C12731_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_29_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_29_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_29_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_29_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_29_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_29_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_29_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_29_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_29_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_29_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_29_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_29_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_29_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_29_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_29_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_29_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_29_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_29_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_29_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_29_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_29_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_29_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_29_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_29_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_29_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_29_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_29_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_29_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_29_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_29_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_29_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_29_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_29_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_29_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_29_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_29_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_29_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_29_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_29_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_29_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_29_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_29_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_29_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_29_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_29_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_29_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_29_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_29_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_29_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_29_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_29_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_29_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_29_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_29_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_29_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_29_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_29_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_29_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_29_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_29_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_29_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_29_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_29_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_29_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N248, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N252, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N254, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N256, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N258, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N260, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N262, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N264, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N266, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N268, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N270, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N272, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N274, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N276, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N278, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N280, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N282, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N284, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N286, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N288, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N290, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N292, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N294, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N296, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N298, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N300, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N302, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N304, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N306, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N308, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N310, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N249, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N251, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N253, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N255, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N257, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N259, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N261, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N263, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N265, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N267, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N269, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N271, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N273, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N275, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N277, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N279, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N281, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N283, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N285, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N287, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N289, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N291, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N293, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N295, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N297, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N299, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N301, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N303, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N305, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N307, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N309, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N311, 
         -- Connections to port 'Z'
         Z(0) => N314 );
   C12732_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_28_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_28_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_28_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_28_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_28_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_28_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_28_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_28_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_28_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_28_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_28_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_28_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_28_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_28_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_28_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_28_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_28_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_28_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_28_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_28_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_28_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_28_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_28_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_28_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_28_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_28_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_28_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_28_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_28_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_28_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_28_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_28_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_28_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_28_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_28_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_28_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_28_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_28_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_28_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_28_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_28_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_28_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_28_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_28_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_28_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_28_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_28_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_28_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_28_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_28_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_28_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_28_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_28_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_28_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_28_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_28_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_28_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_28_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_28_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_28_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_28_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_28_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_28_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_28_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N248, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N252, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N254, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N256, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N258, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N260, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N262, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N264, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N266, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N268, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N270, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N272, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N274, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N276, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N278, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N280, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N282, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N284, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N286, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N288, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N290, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N292, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N294, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N296, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N298, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N300, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N302, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N304, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N306, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N308, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N310, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N249, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N251, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N253, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N255, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N257, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N259, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N261, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N263, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N265, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N267, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N269, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N271, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N273, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N275, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N277, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N279, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N281, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N283, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N285, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N287, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N289, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N291, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N293, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N295, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N297, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N299, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N301, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N303, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N305, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N307, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N309, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N311, 
         -- Connections to port 'Z'
         Z(0) => N315 );
   C12733_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_27_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_27_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_27_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_27_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_27_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_27_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_27_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_27_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_27_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_27_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_27_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_27_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_27_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_27_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_27_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_27_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_27_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_27_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_27_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_27_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_27_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_27_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_27_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_27_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_27_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_27_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_27_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_27_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_27_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_27_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_27_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_27_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_27_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_27_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_27_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_27_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_27_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_27_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_27_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_27_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_27_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_27_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_27_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_27_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_27_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_27_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_27_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_27_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_27_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_27_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_27_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_27_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_27_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_27_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_27_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_27_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_27_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_27_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_27_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_27_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_27_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_27_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_27_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_27_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N248, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N252, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N254, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N256, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N258, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N260, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N262, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N264, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N266, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N268, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N270, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N272, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N274, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N276, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N278, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N280, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N282, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N284, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N286, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N288, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N290, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N292, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N294, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N296, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N298, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N300, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N302, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N304, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N306, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N308, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N310, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N249, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N251, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N253, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N255, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N257, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N259, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N261, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N263, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N265, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N267, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N269, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N271, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N273, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N275, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N277, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N279, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N281, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N283, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N285, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N287, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N289, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N291, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N293, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N295, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N297, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N299, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N301, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N303, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N305, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N307, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N309, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N311, 
         -- Connections to port 'Z'
         Z(0) => N316 );
   C12734_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_26_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_26_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_26_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_26_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_26_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_26_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_26_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_26_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_26_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_26_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_26_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_26_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_26_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_26_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_26_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_26_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_26_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_26_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_26_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_26_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_26_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_26_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_26_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_26_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_26_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_26_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_26_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_26_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_26_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_26_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_26_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_26_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_26_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_26_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_26_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_26_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_26_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_26_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_26_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_26_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_26_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_26_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_26_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_26_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_26_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_26_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_26_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_26_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_26_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_26_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_26_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_26_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_26_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_26_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_26_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_26_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_26_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_26_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_26_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_26_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_26_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_26_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_26_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_26_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N248, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N252, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N254, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N256, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N258, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N260, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N262, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N264, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N266, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N268, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N270, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N272, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N274, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N276, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N278, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N280, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N282, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N284, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N286, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N288, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N290, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N292, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N294, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N296, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N298, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N300, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N302, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N304, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N306, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N308, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N310, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N249, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N251, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N253, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N255, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N257, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N259, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N261, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N263, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N265, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N267, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N269, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N271, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N273, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N275, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N277, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N279, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N281, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N283, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N285, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N287, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N289, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N291, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N293, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N295, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N297, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N299, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N301, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N303, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N305, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N307, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N309, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N311, 
         -- Connections to port 'Z'
         Z(0) => N317 );
   C12735_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_25_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_25_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_25_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_25_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_25_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_25_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_25_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_25_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_25_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_25_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_25_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_25_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_25_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_25_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_25_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_25_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_25_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_25_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_25_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_25_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_25_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_25_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_25_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_25_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_25_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_25_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_25_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_25_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_25_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_25_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_25_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_25_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_25_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_25_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_25_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_25_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_25_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_25_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_25_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_25_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_25_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_25_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_25_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_25_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_25_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_25_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_25_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_25_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_25_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_25_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_25_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_25_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_25_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_25_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_25_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_25_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_25_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_25_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_25_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_25_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_25_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_25_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_25_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_25_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N248, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N252, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N254, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N256, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N258, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N260, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N262, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N264, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N266, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N268, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N270, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N272, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N274, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N276, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N278, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N280, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N282, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N284, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N286, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N288, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N290, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N292, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N294, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N296, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N298, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N300, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N302, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N304, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N306, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N308, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N310, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N249, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N251, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N253, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N255, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N257, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N259, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N261, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N263, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N265, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N267, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N269, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N271, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N273, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N275, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N277, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N279, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N281, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N283, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N285, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N287, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N289, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N291, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N293, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N295, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N297, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N299, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N301, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N303, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N305, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N307, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N309, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N311, 
         -- Connections to port 'Z'
         Z(0) => N318 );
   C12736_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_24_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_24_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_24_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_24_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_24_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_24_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_24_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_24_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_24_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_24_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_24_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_24_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_24_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_24_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_24_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_24_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_24_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_24_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_24_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_24_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_24_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_24_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_24_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_24_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_24_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_24_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_24_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_24_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_24_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_24_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_24_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_24_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_24_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_24_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_24_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_24_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_24_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_24_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_24_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_24_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_24_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_24_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_24_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_24_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_24_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_24_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_24_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_24_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_24_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_24_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_24_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_24_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_24_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_24_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_24_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_24_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_24_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_24_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_24_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_24_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_24_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_24_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_24_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_24_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N248, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N252, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N254, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N256, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N258, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N260, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N262, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N264, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N266, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N268, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N270, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N272, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N274, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N276, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N278, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N280, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N282, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N284, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N286, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N288, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N290, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N292, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N294, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N296, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N298, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N300, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N302, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N304, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N306, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N308, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N310, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N249, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N251, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N253, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N255, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N257, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N259, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N261, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N263, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N265, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N267, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N269, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N271, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N273, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N275, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N277, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N279, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N281, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N283, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N285, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N287, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N289, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N291, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N293, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N295, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N297, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N299, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N301, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N303, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N305, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N307, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N309, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N311, 
         -- Connections to port 'Z'
         Z(0) => N319 );
   C12737_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_23_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_23_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_23_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_23_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_23_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_23_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_23_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_23_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_23_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_23_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_23_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_23_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_23_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_23_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_23_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_23_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_23_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_23_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_23_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_23_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_23_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_23_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_23_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_23_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_23_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_23_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_23_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_23_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_23_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_23_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_23_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_23_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_23_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_23_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_23_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_23_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_23_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_23_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_23_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_23_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_23_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_23_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_23_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_23_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_23_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_23_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_23_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_23_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_23_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_23_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_23_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_23_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_23_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_23_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_23_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_23_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_23_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_23_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_23_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_23_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_23_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_23_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_23_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_23_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N248, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N252, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N254, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N256, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N258, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N260, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N262, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N264, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N266, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N268, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N270, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N272, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N274, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N276, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N278, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N280, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N282, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N284, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N286, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N288, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N290, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N292, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N294, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N296, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N298, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N300, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N302, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N304, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N306, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N308, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N310, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N249, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N251, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N253, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N255, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N257, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N259, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N261, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N263, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N265, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N267, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N269, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N271, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N273, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N275, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N277, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N279, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N281, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N283, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N285, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N287, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N289, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N291, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N293, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N295, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N297, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N299, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N301, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N303, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N305, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N307, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N309, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N311, 
         -- Connections to port 'Z'
         Z(0) => N320 );
   C12738_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_22_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_22_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_22_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_22_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_22_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_22_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_22_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_22_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_22_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_22_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_22_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_22_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_22_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_22_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_22_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_22_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_22_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_22_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_22_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_22_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_22_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_22_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_22_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_22_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_22_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_22_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_22_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_22_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_22_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_22_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_22_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_22_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_22_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_22_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_22_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_22_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_22_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_22_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_22_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_22_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_22_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_22_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_22_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_22_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_22_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_22_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_22_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_22_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_22_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_22_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_22_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_22_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_22_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_22_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_22_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_22_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_22_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_22_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_22_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_22_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_22_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_22_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_22_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_22_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N248, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N252, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N254, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N256, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N258, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N260, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N262, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N264, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N266, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N268, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N270, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N272, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N274, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N276, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N278, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N280, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N282, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N284, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N286, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N288, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N290, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N292, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N294, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N296, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N298, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N300, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N302, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N304, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N306, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N308, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N310, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N249, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N251, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N253, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N255, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N257, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N259, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N261, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N263, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N265, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N267, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N269, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N271, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N273, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N275, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N277, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N279, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N281, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N283, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N285, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N287, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N289, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N291, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N293, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N295, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N297, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N299, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N301, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N303, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N305, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N307, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N309, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N311, 
         -- Connections to port 'Z'
         Z(0) => N321 );
   C12739_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_21_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_21_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_21_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_21_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_21_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_21_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_21_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_21_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_21_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_21_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_21_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_21_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_21_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_21_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_21_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_21_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_21_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_21_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_21_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_21_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_21_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_21_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_21_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_21_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_21_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_21_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_21_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_21_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_21_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_21_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_21_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_21_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_21_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_21_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_21_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_21_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_21_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_21_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_21_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_21_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_21_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_21_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_21_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_21_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_21_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_21_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_21_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_21_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_21_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_21_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_21_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_21_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_21_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_21_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_21_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_21_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_21_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_21_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_21_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_21_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_21_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_21_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_21_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_21_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N248, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N252, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N254, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N256, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N258, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N260, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N262, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N264, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N266, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N268, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N270, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N272, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N274, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N276, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N278, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N280, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N282, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N284, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N286, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N288, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N290, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N292, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N294, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N296, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N298, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N300, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N302, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N304, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N306, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N308, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N310, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N249, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N251, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N253, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N255, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N257, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N259, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N261, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N263, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N265, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N267, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N269, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N271, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N273, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N275, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N277, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N279, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N281, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N283, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N285, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N287, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N289, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N291, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N293, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N295, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N297, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N299, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N301, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N303, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N305, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N307, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N309, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N311, 
         -- Connections to port 'Z'
         Z(0) => N322 );
   C12740_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_20_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_20_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_20_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_20_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_20_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_20_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_20_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_20_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_20_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_20_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_20_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_20_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_20_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_20_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_20_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_20_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_20_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_20_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_20_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_20_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_20_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_20_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_20_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_20_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_20_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_20_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_20_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_20_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_20_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_20_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_20_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_20_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_20_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_20_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_20_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_20_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_20_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_20_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_20_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_20_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_20_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_20_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_20_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_20_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_20_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_20_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_20_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_20_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_20_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_20_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_20_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_20_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_20_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_20_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_20_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_20_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_20_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_20_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_20_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_20_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_20_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_20_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_20_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_20_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N248, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N252, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N254, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N256, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N258, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N260, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N262, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N264, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N266, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N268, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N270, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N272, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N274, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N276, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N278, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N280, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N282, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N284, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N286, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N288, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N290, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N292, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N294, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N296, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N298, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N300, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N302, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N304, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N306, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N308, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N310, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N249, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N251, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N253, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N255, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N257, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N259, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N261, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N263, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N265, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N267, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N269, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N271, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N273, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N275, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N277, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N279, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N281, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N283, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N285, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N287, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N289, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N291, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N293, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N295, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N297, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N299, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N301, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N303, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N305, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N307, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N309, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N311, 
         -- Connections to port 'Z'
         Z(0) => N323 );
   C12741_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_19_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_19_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_19_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_19_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_19_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_19_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_19_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_19_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_19_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_19_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_19_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_19_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_19_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_19_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_19_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_19_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_19_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_19_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_19_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_19_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_19_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_19_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_19_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_19_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_19_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_19_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_19_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_19_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_19_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_19_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_19_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_19_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_19_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_19_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_19_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_19_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_19_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_19_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_19_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_19_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_19_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_19_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_19_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_19_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_19_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_19_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_19_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_19_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_19_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_19_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_19_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_19_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_19_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_19_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_19_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_19_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_19_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_19_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_19_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_19_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_19_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_19_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_19_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_19_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N248, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N252, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N254, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N256, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N258, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N260, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N262, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N264, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N266, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N268, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N270, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N272, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N274, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N276, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N278, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N280, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N282, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N284, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N286, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N288, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N290, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N292, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N294, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N296, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N298, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N300, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N302, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N304, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N306, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N308, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N310, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N249, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N251, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N253, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N255, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N257, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N259, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N261, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N263, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N265, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N267, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N269, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N271, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N273, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N275, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N277, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N279, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N281, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N283, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N285, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N287, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N289, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N291, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N293, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N295, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N297, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N299, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N301, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N303, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N305, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N307, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N309, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N311, 
         -- Connections to port 'Z'
         Z(0) => N324 );
   C12742_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_18_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_18_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_18_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_18_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_18_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_18_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_18_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_18_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_18_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_18_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_18_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_18_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_18_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_18_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_18_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_18_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_18_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_18_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_18_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_18_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_18_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_18_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_18_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_18_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_18_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_18_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_18_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_18_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_18_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_18_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_18_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_18_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_18_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_18_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_18_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_18_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_18_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_18_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_18_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_18_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_18_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_18_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_18_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_18_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_18_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_18_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_18_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_18_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_18_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_18_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_18_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_18_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_18_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_18_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_18_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_18_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_18_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_18_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_18_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_18_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_18_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_18_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_18_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_18_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N248, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N252, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N254, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N256, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N258, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N260, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N262, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N264, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N266, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N268, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N270, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N272, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N274, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N276, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N278, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N280, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N282, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N284, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N286, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N288, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N290, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N292, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N294, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N296, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N298, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N300, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N302, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N304, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N306, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N308, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N310, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N249, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N251, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N253, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N255, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N257, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N259, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N261, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N263, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N265, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N267, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N269, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N271, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N273, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N275, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N277, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N279, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N281, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N283, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N285, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N287, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N289, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N291, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N293, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N295, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N297, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N299, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N301, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N303, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N305, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N307, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N309, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N311, 
         -- Connections to port 'Z'
         Z(0) => N325 );
   C12743_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_17_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_17_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_17_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_17_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_17_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_17_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_17_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_17_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_17_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_17_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_17_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_17_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_17_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_17_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_17_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_17_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_17_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_17_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_17_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_17_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_17_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_17_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_17_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_17_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_17_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_17_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_17_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_17_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_17_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_17_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_17_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_17_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_17_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_17_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_17_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_17_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_17_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_17_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_17_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_17_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_17_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_17_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_17_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_17_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_17_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_17_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_17_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_17_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_17_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_17_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_17_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_17_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_17_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_17_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_17_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_17_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_17_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_17_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_17_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_17_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_17_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_17_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_17_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_17_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N248, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N252, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N254, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N256, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N258, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N260, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N262, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N264, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N266, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N268, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N270, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N272, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N274, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N276, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N278, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N280, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N282, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N284, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N286, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N288, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N290, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N292, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N294, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N296, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N298, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N300, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N302, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N304, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N306, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N308, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N310, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N249, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N251, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N253, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N255, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N257, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N259, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N261, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N263, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N265, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N267, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N269, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N271, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N273, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N275, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N277, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N279, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N281, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N283, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N285, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N287, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N289, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N291, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N293, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N295, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N297, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N299, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N301, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N303, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N305, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N307, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N309, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N311, 
         -- Connections to port 'Z'
         Z(0) => N326 );
   C12744_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_16_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_16_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_16_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_16_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_16_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_16_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_16_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_16_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_16_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_16_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_16_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_16_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_16_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_16_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_16_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_16_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_16_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_16_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_16_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_16_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_16_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_16_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_16_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_16_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_16_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_16_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_16_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_16_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_16_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_16_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_16_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_16_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_16_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_16_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_16_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_16_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_16_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_16_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_16_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_16_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_16_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_16_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_16_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_16_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_16_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_16_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_16_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_16_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_16_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_16_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_16_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_16_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_16_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_16_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_16_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_16_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_16_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_16_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_16_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_16_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_16_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_16_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_16_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_16_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N248, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N252, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N254, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N256, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N258, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N260, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N262, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N264, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N266, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N268, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N270, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N272, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N274, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N276, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N278, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N280, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N282, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N284, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N286, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N288, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N290, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N292, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N294, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N296, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N298, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N300, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N302, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N304, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N306, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N308, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N310, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N249, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N251, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N253, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N255, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N257, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N259, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N261, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N263, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N265, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N267, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N269, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N271, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N273, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N275, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N277, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N279, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N281, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N283, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N285, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N287, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N289, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N291, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N293, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N295, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N297, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N299, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N301, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N303, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N305, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N307, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N309, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N311, 
         -- Connections to port 'Z'
         Z(0) => N327 );
   C12745_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_15_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_15_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_15_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_15_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_15_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_15_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_15_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_15_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_15_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_15_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_15_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_15_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_15_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_15_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_15_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_15_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_15_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_15_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_15_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_15_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_15_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_15_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_15_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_15_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_15_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_15_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_15_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_15_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_15_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_15_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_15_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_15_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_15_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_15_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_15_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_15_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_15_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_15_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_15_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_15_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_15_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_15_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_15_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_15_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_15_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_15_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_15_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_15_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_15_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_15_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_15_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_15_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_15_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_15_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_15_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_15_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_15_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_15_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_15_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_15_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_15_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_15_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_15_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_15_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N248, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N252, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N254, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N256, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N258, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N260, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N262, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N264, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N266, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N268, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N270, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N272, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N274, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N276, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N278, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N280, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N282, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N284, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N286, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N288, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N290, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N292, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N294, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N296, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N298, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N300, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N302, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N304, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N306, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N308, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N310, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N249, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N251, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N253, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N255, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N257, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N259, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N261, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N263, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N265, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N267, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N269, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N271, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N273, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N275, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N277, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N279, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N281, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N283, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N285, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N287, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N289, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N291, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N293, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N295, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N297, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N299, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N301, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N303, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N305, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N307, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N309, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N311, 
         -- Connections to port 'Z'
         Z(0) => N328 );
   C12746_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_14_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_14_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_14_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_14_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_14_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_14_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_14_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_14_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_14_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_14_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_14_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_14_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_14_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_14_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_14_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_14_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_14_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_14_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_14_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_14_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_14_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_14_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_14_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_14_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_14_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_14_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_14_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_14_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_14_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_14_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_14_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_14_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_14_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_14_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_14_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_14_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_14_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_14_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_14_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_14_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_14_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_14_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_14_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_14_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_14_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_14_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_14_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_14_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_14_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_14_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_14_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_14_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_14_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_14_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_14_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_14_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_14_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_14_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_14_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_14_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_14_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_14_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_14_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_14_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N248, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N252, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N254, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N256, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N258, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N260, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N262, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N264, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N266, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N268, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N270, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N272, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N274, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N276, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N278, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N280, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N282, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N284, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N286, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N288, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N290, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N292, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N294, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N296, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N298, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N300, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N302, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N304, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N306, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N308, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N310, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N249, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N251, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N253, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N255, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N257, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N259, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N261, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N263, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N265, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N267, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N269, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N271, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N273, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N275, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N277, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N279, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N281, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N283, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N285, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N287, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N289, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N291, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N293, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N295, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N297, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N299, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N301, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N303, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N305, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N307, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N309, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N311, 
         -- Connections to port 'Z'
         Z(0) => N329 );
   C12747_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_13_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_13_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_13_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_13_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_13_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_13_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_13_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_13_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_13_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_13_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_13_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_13_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_13_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_13_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_13_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_13_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_13_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_13_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_13_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_13_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_13_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_13_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_13_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_13_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_13_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_13_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_13_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_13_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_13_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_13_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_13_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_13_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_13_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_13_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_13_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_13_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_13_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_13_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_13_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_13_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_13_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_13_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_13_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_13_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_13_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_13_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_13_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_13_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_13_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_13_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_13_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_13_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_13_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_13_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_13_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_13_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_13_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_13_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_13_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_13_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_13_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_13_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_13_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_13_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N248, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N252, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N254, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N256, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N258, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N260, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N262, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N264, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N266, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N268, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N270, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N272, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N274, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N276, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N278, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N280, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N282, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N284, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N286, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N288, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N290, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N292, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N294, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N296, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N298, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N300, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N302, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N304, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N306, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N308, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N310, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N249, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N251, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N253, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N255, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N257, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N259, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N261, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N263, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N265, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N267, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N269, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N271, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N273, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N275, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N277, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N279, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N281, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N283, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N285, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N287, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N289, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N291, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N293, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N295, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N297, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N299, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N301, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N303, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N305, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N307, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N309, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N311, 
         -- Connections to port 'Z'
         Z(0) => N330 );
   C12748_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_12_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_12_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_12_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_12_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_12_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_12_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_12_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_12_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_12_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_12_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_12_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_12_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_12_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_12_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_12_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_12_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_12_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_12_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_12_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_12_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_12_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_12_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_12_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_12_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_12_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_12_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_12_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_12_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_12_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_12_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_12_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_12_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_12_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_12_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_12_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_12_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_12_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_12_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_12_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_12_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_12_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_12_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_12_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_12_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_12_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_12_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_12_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_12_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_12_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_12_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_12_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_12_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_12_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_12_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_12_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_12_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_12_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_12_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_12_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_12_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_12_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_12_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_12_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_12_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N248, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N252, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N254, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N256, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N258, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N260, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N262, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N264, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N266, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N268, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N270, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N272, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N274, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N276, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N278, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N280, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N282, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N284, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N286, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N288, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N290, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N292, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N294, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N296, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N298, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N300, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N302, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N304, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N306, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N308, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N310, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N249, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N251, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N253, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N255, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N257, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N259, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N261, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N263, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N265, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N267, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N269, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N271, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N273, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N275, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N277, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N279, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N281, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N283, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N285, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N287, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N289, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N291, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N293, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N295, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N297, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N299, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N301, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N303, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N305, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N307, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N309, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N311, 
         -- Connections to port 'Z'
         Z(0) => N331 );
   C12749_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_11_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_11_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_11_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_11_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_11_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_11_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_11_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_11_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_11_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_11_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_11_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_11_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_11_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_11_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_11_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_11_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_11_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_11_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_11_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_11_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_11_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_11_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_11_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_11_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_11_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_11_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_11_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_11_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_11_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_11_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_11_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_11_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_11_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_11_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_11_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_11_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_11_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_11_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_11_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_11_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_11_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_11_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_11_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_11_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_11_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_11_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_11_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_11_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_11_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_11_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_11_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_11_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_11_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_11_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_11_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_11_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_11_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_11_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_11_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_11_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_11_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_11_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_11_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_11_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N248, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N252, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N254, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N256, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N258, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N260, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N262, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N264, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N266, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N268, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N270, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N272, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N274, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N276, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N278, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N280, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N282, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N284, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N286, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N288, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N290, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N292, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N294, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N296, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N298, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N300, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N302, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N304, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N306, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N308, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N310, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N249, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N251, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N253, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N255, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N257, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N259, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N261, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N263, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N265, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N267, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N269, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N271, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N273, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N275, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N277, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N279, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N281, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N283, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N285, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N287, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N289, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N291, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N293, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N295, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N297, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N299, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N301, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N303, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N305, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N307, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N309, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N311, 
         -- Connections to port 'Z'
         Z(0) => N332 );
   C12750_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_10_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_10_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_10_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_10_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_10_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_10_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_10_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_10_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_10_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_10_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_10_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_10_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_10_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_10_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_10_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_10_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_10_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_10_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_10_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_10_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_10_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_10_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_10_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_10_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_10_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_10_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_10_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_10_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_10_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_10_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_10_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_10_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_10_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_10_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_10_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_10_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_10_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_10_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_10_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_10_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_10_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_10_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_10_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_10_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_10_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_10_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_10_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_10_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_10_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_10_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_10_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_10_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_10_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_10_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_10_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_10_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_10_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_10_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_10_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_10_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_10_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_10_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_10_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_10_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N248, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N252, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N254, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N256, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N258, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N260, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N262, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N264, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N266, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N268, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N270, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N272, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N274, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N276, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N278, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N280, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N282, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N284, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N286, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N288, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N290, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N292, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N294, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N296, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N298, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N300, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N302, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N304, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N306, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N308, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N310, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N249, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N251, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N253, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N255, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N257, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N259, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N261, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N263, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N265, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N267, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N269, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N271, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N273, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N275, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N277, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N279, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N281, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N283, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N285, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N287, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N289, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N291, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N293, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N295, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N297, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N299, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N301, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N303, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N305, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N307, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N309, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N311, 
         -- Connections to port 'Z'
         Z(0) => N333 );
   C12751_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_9_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_9_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_9_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_9_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_9_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_9_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_9_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_9_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_9_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_9_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_9_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_9_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_9_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_9_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_9_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_9_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_9_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_9_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_9_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_9_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_9_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_9_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_9_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_9_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_9_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_9_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_9_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_9_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_9_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_9_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_9_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_9_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_9_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_9_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_9_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_9_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_9_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_9_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_9_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_9_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_9_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_9_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_9_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_9_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_9_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_9_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_9_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_9_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_9_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_9_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_9_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_9_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_9_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_9_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_9_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_9_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_9_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_9_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_9_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_9_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_9_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_9_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_9_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_9_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N248, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N252, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N254, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N256, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N258, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N260, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N262, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N264, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N266, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N268, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N270, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N272, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N274, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N276, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N278, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N280, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N282, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N284, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N286, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N288, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N290, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N292, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N294, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N296, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N298, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N300, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N302, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N304, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N306, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N308, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N310, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N249, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N251, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N253, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N255, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N257, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N259, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N261, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N263, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N265, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N267, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N269, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N271, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N273, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N275, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N277, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N279, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N281, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N283, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N285, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N287, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N289, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N291, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N293, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N295, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N297, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N299, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N301, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N303, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N305, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N307, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N309, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N311, 
         -- Connections to port 'Z'
         Z(0) => N334 );
   C12752_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_8_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_8_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_8_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_8_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_8_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_8_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_8_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_8_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_8_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_8_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_8_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_8_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_8_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_8_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_8_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_8_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_8_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_8_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_8_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_8_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_8_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_8_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_8_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_8_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_8_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_8_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_8_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_8_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_8_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_8_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_8_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_8_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_8_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_8_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_8_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_8_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_8_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_8_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_8_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_8_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_8_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_8_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_8_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_8_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_8_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_8_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_8_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_8_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_8_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_8_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_8_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_8_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_8_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_8_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_8_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_8_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_8_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_8_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_8_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_8_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_8_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_8_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_8_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_8_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N248, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N252, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N254, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N256, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N258, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N260, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N262, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N264, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N266, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N268, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N270, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N272, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N274, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N276, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N278, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N280, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N282, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N284, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N286, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N288, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N290, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N292, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N294, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N296, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N298, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N300, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N302, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N304, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N306, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N308, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N310, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N249, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N251, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N253, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N255, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N257, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N259, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N261, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N263, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N265, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N267, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N269, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N271, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N273, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N275, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N277, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N279, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N281, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N283, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N285, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N287, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N289, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N291, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N293, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N295, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N297, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N299, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N301, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N303, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N305, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N307, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N309, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N311, 
         -- Connections to port 'Z'
         Z(0) => N335 );
   C12753_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_7_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_7_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_7_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_7_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_7_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_7_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_7_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_7_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_7_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_7_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_7_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_7_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_7_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_7_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_7_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_7_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_7_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_7_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_7_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_7_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_7_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_7_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_7_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_7_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_7_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_7_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_7_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_7_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_7_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_7_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_7_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_7_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_7_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_7_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_7_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_7_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_7_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_7_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_7_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_7_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_7_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_7_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_7_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_7_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_7_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_7_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_7_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_7_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_7_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_7_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_7_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_7_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_7_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_7_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_7_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_7_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_7_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_7_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_7_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_7_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_7_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_7_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_7_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_7_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N248, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N252, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N254, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N256, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N258, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N260, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N262, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N264, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N266, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N268, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N270, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N272, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N274, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N276, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N278, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N280, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N282, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N284, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N286, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N288, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N290, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N292, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N294, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N296, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N298, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N300, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N302, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N304, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N306, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N308, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N310, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N249, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N251, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N253, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N255, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N257, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N259, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N261, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N263, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N265, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N267, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N269, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N271, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N273, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N275, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N277, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N279, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N281, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N283, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N285, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N287, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N289, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N291, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N293, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N295, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N297, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N299, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N301, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N303, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N305, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N307, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N309, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N311, 
         -- Connections to port 'Z'
         Z(0) => N336 );
   C12754_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_6_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_6_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_6_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_6_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_6_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_6_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_6_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_6_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_6_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_6_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_6_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_6_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_6_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_6_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_6_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_6_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_6_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_6_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_6_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_6_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_6_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_6_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_6_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_6_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_6_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_6_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_6_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_6_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_6_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_6_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_6_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_6_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_6_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_6_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_6_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_6_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_6_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_6_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_6_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_6_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_6_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_6_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_6_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_6_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_6_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_6_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_6_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_6_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_6_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_6_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_6_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_6_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_6_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_6_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_6_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_6_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_6_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_6_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_6_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_6_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_6_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_6_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_6_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_6_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N248, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N252, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N254, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N256, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N258, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N260, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N262, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N264, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N266, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N268, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N270, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N272, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N274, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N276, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N278, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N280, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N282, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N284, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N286, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N288, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N290, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N292, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N294, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N296, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N298, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N300, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N302, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N304, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N306, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N308, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N310, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N249, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N251, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N253, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N255, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N257, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N259, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N261, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N263, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N265, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N267, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N269, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N271, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N273, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N275, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N277, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N279, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N281, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N283, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N285, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N287, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N289, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N291, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N293, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N295, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N297, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N299, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N301, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N303, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N305, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N307, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N309, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N311, 
         -- Connections to port 'Z'
         Z(0) => N337 );
   C12755_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_5_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_5_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_5_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_5_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_5_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_5_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_5_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_5_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_5_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_5_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_5_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_5_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_5_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_5_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_5_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_5_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_5_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_5_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_5_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_5_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_5_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_5_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_5_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_5_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_5_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_5_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_5_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_5_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_5_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_5_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_5_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_5_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_5_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_5_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_5_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_5_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_5_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_5_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_5_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_5_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_5_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_5_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_5_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_5_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_5_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_5_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_5_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_5_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_5_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_5_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_5_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_5_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_5_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_5_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_5_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_5_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_5_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_5_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_5_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_5_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_5_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_5_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_5_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_5_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N248, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N252, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N254, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N256, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N258, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N260, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N262, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N264, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N266, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N268, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N270, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N272, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N274, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N276, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N278, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N280, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N282, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N284, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N286, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N288, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N290, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N292, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N294, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N296, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N298, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N300, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N302, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N304, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N306, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N308, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N310, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N249, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N251, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N253, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N255, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N257, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N259, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N261, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N263, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N265, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N267, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N269, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N271, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N273, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N275, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N277, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N279, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N281, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N283, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N285, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N287, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N289, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N291, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N293, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N295, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N297, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N299, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N301, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N303, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N305, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N307, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N309, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N311, 
         -- Connections to port 'Z'
         Z(0) => N338 );
   C12756_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_4_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_4_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_4_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_4_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_4_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_4_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_4_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_4_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_4_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_4_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_4_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_4_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_4_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_4_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_4_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_4_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_4_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_4_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_4_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_4_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_4_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_4_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_4_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_4_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_4_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_4_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_4_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_4_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_4_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_4_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_4_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_4_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_4_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_4_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_4_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_4_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_4_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_4_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_4_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_4_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_4_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_4_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_4_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_4_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_4_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_4_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_4_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_4_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_4_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_4_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_4_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_4_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_4_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_4_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_4_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_4_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_4_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_4_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_4_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_4_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_4_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_4_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_4_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_4_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N248, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N252, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N254, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N256, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N258, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N260, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N262, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N264, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N266, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N268, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N270, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N272, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N274, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N276, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N278, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N280, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N282, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N284, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N286, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N288, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N290, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N292, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N294, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N296, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N298, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N300, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N302, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N304, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N306, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N308, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N310, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N249, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N251, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N253, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N255, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N257, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N259, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N261, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N263, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N265, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N267, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N269, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N271, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N273, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N275, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N277, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N279, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N281, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N283, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N285, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N287, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N289, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N291, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N293, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N295, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N297, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N299, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N301, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N303, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N305, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N307, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N309, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N311, 
         -- Connections to port 'Z'
         Z(0) => N339 );
   C12757_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_3_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_3_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_3_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_3_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_3_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_3_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_3_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_3_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_3_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_3_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_3_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_3_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_3_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_3_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_3_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_3_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_3_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_3_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_3_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_3_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_3_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_3_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_3_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_3_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_3_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_3_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_3_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_3_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_3_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_3_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_3_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_3_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_3_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_3_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_3_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_3_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_3_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_3_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_3_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_3_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_3_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_3_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_3_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_3_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_3_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_3_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_3_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_3_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_3_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_3_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_3_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_3_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_3_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_3_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_3_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_3_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_3_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_3_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_3_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_3_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_3_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_3_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_3_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_3_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N248, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N252, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N254, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N256, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N258, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N260, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N262, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N264, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N266, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N268, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N270, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N272, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N274, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N276, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N278, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N280, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N282, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N284, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N286, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N288, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N290, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N292, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N294, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N296, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N298, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N300, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N302, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N304, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N306, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N308, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N310, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N249, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N251, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N253, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N255, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N257, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N259, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N261, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N263, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N265, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N267, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N269, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N271, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N273, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N275, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N277, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N279, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N281, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N283, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N285, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N287, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N289, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N291, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N293, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N295, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N297, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N299, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N301, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N303, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N305, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N307, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N309, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N311, 
         -- Connections to port 'Z'
         Z(0) => N340 );
   C12758_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_2_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_2_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_2_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_2_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_2_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_2_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_2_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_2_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_2_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_2_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_2_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_2_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_2_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_2_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_2_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_2_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_2_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_2_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_2_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_2_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_2_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_2_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_2_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_2_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_2_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_2_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_2_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_2_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_2_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_2_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_2_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_2_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_2_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_2_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_2_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_2_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_2_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_2_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_2_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_2_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_2_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_2_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_2_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_2_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_2_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_2_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_2_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_2_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_2_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_2_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_2_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_2_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_2_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_2_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_2_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_2_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_2_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_2_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_2_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_2_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_2_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_2_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_2_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_2_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N248, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N252, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N254, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N256, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N258, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N260, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N262, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N264, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N266, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N268, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N270, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N272, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N274, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N276, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N278, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N280, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N282, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N284, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N286, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N288, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N290, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N292, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N294, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N296, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N298, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N300, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N302, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N304, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N306, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N308, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N310, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N249, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N251, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N253, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N255, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N257, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N259, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N261, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N263, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N265, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N267, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N269, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N271, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N273, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N275, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N277, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N279, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N281, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N283, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N285, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N287, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N289, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N291, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N293, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N295, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N297, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N299, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N301, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N303, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N305, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N307, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N309, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N311, 
         -- Connections to port 'Z'
         Z(0) => N341 );
   C12759_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_1_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_1_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_1_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_1_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_1_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_1_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_1_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_1_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_1_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_1_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_1_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_1_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_1_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_1_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_1_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_1_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_1_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_1_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_1_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_1_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_1_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_1_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_1_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_1_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_1_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_1_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_1_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_1_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_1_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_1_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_1_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_1_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_1_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_1_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_1_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_1_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_1_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_1_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_1_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_1_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_1_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_1_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_1_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_1_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_1_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_1_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_1_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_1_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_1_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_1_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_1_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_1_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_1_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_1_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_1_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_1_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_1_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_1_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_1_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_1_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_1_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_1_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_1_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_1_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N248, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N252, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N254, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N256, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N258, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N260, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N262, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N264, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N266, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N268, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N270, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N272, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N274, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N276, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N278, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N280, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N282, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N284, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N286, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N288, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N290, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N292, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N294, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N296, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N298, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N300, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N302, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N304, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N306, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N308, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N310, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N249, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N251, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N253, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N255, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N257, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N259, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N261, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N263, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N265, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N267, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N269, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N271, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N273, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N275, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N277, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N279, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N281, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N283, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N285, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N287, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N289, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N291, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N293, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N295, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N297, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N299, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N301, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N303, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N305, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N307, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N309, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N311, 
         -- Connections to port 'Z'
         Z(0) => N342 );
   C12760_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_0_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_0_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_0_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_0_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_0_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_0_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_0_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_0_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_0_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_0_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_0_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_0_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_0_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_0_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_0_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_0_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_0_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_0_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_0_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_0_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_0_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_0_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_0_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_0_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_0_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_0_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_0_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_0_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_0_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_0_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_0_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_0_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_0_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_0_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_0_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_0_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_0_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_0_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_0_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_0_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_0_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_0_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_0_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_0_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_0_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_0_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_0_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_0_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_0_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_0_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_0_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_0_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_0_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_0_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_0_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_0_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_0_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_0_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_0_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_0_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_0_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_0_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N248, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N252, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N254, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N256, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N258, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N260, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N262, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N264, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N266, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N268, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N270, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N272, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N274, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N276, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N278, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N280, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N282, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N284, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N286, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N288, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N290, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N292, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N294, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N296, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N298, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N300, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N302, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N304, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N306, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N308, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N310, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N249, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N251, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N253, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N255, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N257, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N259, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N261, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N263, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N265, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N267, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N269, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N271, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N273, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N275, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N277, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N279, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N281, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N283, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N285, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N287, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N289, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N291, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N293, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N295, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N297, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N299, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N301, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N303, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N305, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N307, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N309, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N311, 
         -- Connections to port 'Z'
         Z(0) => N343 );
   C12891_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_31_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_31_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_31_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_31_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_31_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_31_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_31_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_31_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_31_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_31_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_31_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_31_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_31_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_31_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_31_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_31_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_31_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_31_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_31_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_31_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_31_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_31_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_31_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_31_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_31_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_31_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_31_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_31_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_31_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_31_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_31_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_31_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_31_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_31_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_31_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_31_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_31_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_31_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_31_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_31_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_31_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_31_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_31_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_31_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_31_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_31_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_31_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_31_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_31_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_31_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_31_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_31_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_31_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_31_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_31_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_31_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_31_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_31_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_31_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_31_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_31_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_31_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_31_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_31_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N410, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N412, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N414, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N416, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N418, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N420, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N422, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N424, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N426, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N428, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N430, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N432, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N434, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N436, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N438, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N440, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N442, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N444, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N446, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N448, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N450, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N452, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N454, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N456, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N458, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N460, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N462, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N464, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N466, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N468, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N470, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N472, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N411, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N413, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N415, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N417, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N419, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N421, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N423, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N425, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N427, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N429, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N431, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N433, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N435, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N437, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N439, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N441, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N443, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N445, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N447, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N449, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N451, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N453, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N455, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N457, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N459, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N461, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N463, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N465, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N467, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N469, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N471, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N473, 
         -- Connections to port 'Z'
         Z(0) => N474 );
   C12892_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_30_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_30_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_30_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_30_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_30_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_30_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_30_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_30_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_30_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_30_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_30_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_30_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_30_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_30_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_30_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_30_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_30_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_30_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_30_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_30_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_30_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_30_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_30_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_30_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_30_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_30_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_30_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_30_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_30_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_30_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_30_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_30_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_30_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_30_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_30_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_30_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_30_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_30_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_30_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_30_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_30_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_30_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_30_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_30_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_30_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_30_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_30_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_30_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_30_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_30_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_30_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_30_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_30_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_30_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_30_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_30_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_30_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_30_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_30_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_30_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_30_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_30_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_30_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_30_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N410, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N412, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N414, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N416, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N418, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N420, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N422, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N424, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N426, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N428, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N430, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N432, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N434, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N436, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N438, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N440, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N442, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N444, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N446, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N448, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N450, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N452, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N454, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N456, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N458, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N460, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N462, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N464, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N466, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N468, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N470, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N472, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N411, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N413, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N415, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N417, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N419, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N421, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N423, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N425, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N427, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N429, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N431, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N433, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N435, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N437, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N439, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N441, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N443, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N445, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N447, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N449, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N451, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N453, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N455, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N457, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N459, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N461, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N463, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N465, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N467, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N469, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N471, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N473, 
         -- Connections to port 'Z'
         Z(0) => N475 );
   C12893_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_29_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_29_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_29_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_29_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_29_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_29_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_29_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_29_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_29_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_29_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_29_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_29_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_29_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_29_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_29_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_29_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_29_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_29_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_29_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_29_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_29_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_29_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_29_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_29_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_29_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_29_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_29_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_29_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_29_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_29_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_29_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_29_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_29_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_29_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_29_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_29_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_29_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_29_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_29_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_29_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_29_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_29_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_29_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_29_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_29_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_29_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_29_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_29_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_29_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_29_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_29_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_29_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_29_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_29_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_29_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_29_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_29_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_29_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_29_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_29_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_29_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_29_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_29_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_29_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N410, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N412, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N414, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N416, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N418, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N420, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N422, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N424, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N426, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N428, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N430, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N432, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N434, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N436, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N438, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N440, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N442, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N444, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N446, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N448, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N450, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N452, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N454, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N456, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N458, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N460, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N462, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N464, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N466, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N468, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N470, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N472, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N411, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N413, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N415, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N417, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N419, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N421, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N423, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N425, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N427, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N429, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N431, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N433, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N435, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N437, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N439, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N441, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N443, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N445, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N447, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N449, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N451, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N453, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N455, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N457, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N459, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N461, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N463, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N465, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N467, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N469, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N471, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N473, 
         -- Connections to port 'Z'
         Z(0) => N476 );
   C12894_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_28_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_28_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_28_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_28_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_28_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_28_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_28_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_28_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_28_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_28_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_28_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_28_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_28_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_28_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_28_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_28_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_28_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_28_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_28_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_28_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_28_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_28_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_28_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_28_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_28_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_28_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_28_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_28_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_28_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_28_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_28_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_28_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_28_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_28_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_28_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_28_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_28_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_28_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_28_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_28_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_28_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_28_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_28_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_28_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_28_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_28_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_28_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_28_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_28_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_28_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_28_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_28_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_28_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_28_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_28_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_28_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_28_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_28_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_28_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_28_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_28_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_28_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_28_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_28_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N410, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N412, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N414, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N416, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N418, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N420, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N422, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N424, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N426, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N428, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N430, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N432, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N434, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N436, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N438, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N440, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N442, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N444, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N446, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N448, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N450, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N452, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N454, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N456, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N458, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N460, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N462, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N464, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N466, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N468, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N470, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N472, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N411, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N413, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N415, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N417, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N419, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N421, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N423, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N425, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N427, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N429, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N431, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N433, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N435, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N437, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N439, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N441, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N443, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N445, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N447, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N449, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N451, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N453, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N455, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N457, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N459, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N461, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N463, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N465, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N467, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N469, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N471, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N473, 
         -- Connections to port 'Z'
         Z(0) => N477 );
   C12895_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_27_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_27_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_27_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_27_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_27_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_27_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_27_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_27_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_27_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_27_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_27_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_27_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_27_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_27_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_27_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_27_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_27_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_27_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_27_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_27_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_27_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_27_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_27_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_27_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_27_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_27_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_27_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_27_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_27_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_27_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_27_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_27_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_27_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_27_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_27_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_27_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_27_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_27_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_27_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_27_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_27_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_27_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_27_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_27_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_27_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_27_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_27_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_27_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_27_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_27_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_27_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_27_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_27_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_27_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_27_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_27_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_27_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_27_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_27_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_27_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_27_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_27_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_27_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_27_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N410, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N412, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N414, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N416, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N418, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N420, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N422, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N424, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N426, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N428, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N430, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N432, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N434, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N436, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N438, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N440, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N442, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N444, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N446, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N448, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N450, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N452, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N454, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N456, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N458, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N460, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N462, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N464, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N466, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N468, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N470, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N472, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N411, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N413, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N415, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N417, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N419, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N421, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N423, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N425, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N427, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N429, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N431, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N433, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N435, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N437, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N439, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N441, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N443, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N445, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N447, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N449, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N451, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N453, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N455, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N457, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N459, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N461, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N463, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N465, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N467, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N469, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N471, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N473, 
         -- Connections to port 'Z'
         Z(0) => N478 );
   C12896_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_26_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_26_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_26_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_26_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_26_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_26_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_26_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_26_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_26_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_26_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_26_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_26_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_26_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_26_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_26_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_26_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_26_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_26_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_26_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_26_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_26_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_26_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_26_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_26_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_26_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_26_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_26_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_26_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_26_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_26_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_26_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_26_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_26_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_26_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_26_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_26_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_26_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_26_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_26_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_26_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_26_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_26_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_26_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_26_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_26_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_26_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_26_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_26_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_26_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_26_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_26_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_26_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_26_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_26_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_26_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_26_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_26_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_26_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_26_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_26_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_26_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_26_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_26_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_26_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N410, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N412, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N414, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N416, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N418, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N420, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N422, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N424, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N426, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N428, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N430, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N432, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N434, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N436, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N438, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N440, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N442, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N444, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N446, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N448, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N450, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N452, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N454, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N456, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N458, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N460, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N462, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N464, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N466, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N468, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N470, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N472, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N411, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N413, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N415, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N417, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N419, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N421, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N423, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N425, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N427, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N429, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N431, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N433, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N435, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N437, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N439, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N441, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N443, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N445, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N447, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N449, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N451, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N453, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N455, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N457, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N459, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N461, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N463, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N465, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N467, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N469, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N471, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N473, 
         -- Connections to port 'Z'
         Z(0) => N479 );
   C12897_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_25_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_25_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_25_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_25_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_25_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_25_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_25_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_25_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_25_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_25_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_25_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_25_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_25_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_25_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_25_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_25_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_25_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_25_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_25_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_25_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_25_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_25_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_25_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_25_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_25_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_25_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_25_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_25_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_25_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_25_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_25_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_25_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_25_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_25_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_25_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_25_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_25_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_25_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_25_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_25_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_25_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_25_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_25_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_25_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_25_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_25_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_25_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_25_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_25_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_25_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_25_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_25_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_25_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_25_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_25_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_25_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_25_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_25_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_25_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_25_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_25_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_25_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_25_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_25_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N410, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N412, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N414, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N416, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N418, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N420, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N422, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N424, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N426, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N428, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N430, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N432, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N434, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N436, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N438, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N440, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N442, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N444, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N446, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N448, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N450, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N452, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N454, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N456, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N458, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N460, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N462, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N464, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N466, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N468, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N470, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N472, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N411, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N413, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N415, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N417, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N419, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N421, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N423, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N425, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N427, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N429, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N431, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N433, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N435, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N437, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N439, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N441, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N443, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N445, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N447, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N449, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N451, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N453, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N455, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N457, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N459, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N461, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N463, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N465, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N467, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N469, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N471, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N473, 
         -- Connections to port 'Z'
         Z(0) => N480 );
   C12898_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_24_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_24_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_24_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_24_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_24_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_24_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_24_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_24_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_24_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_24_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_24_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_24_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_24_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_24_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_24_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_24_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_24_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_24_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_24_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_24_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_24_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_24_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_24_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_24_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_24_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_24_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_24_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_24_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_24_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_24_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_24_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_24_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_24_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_24_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_24_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_24_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_24_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_24_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_24_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_24_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_24_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_24_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_24_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_24_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_24_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_24_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_24_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_24_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_24_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_24_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_24_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_24_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_24_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_24_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_24_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_24_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_24_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_24_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_24_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_24_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_24_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_24_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_24_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_24_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N410, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N412, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N414, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N416, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N418, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N420, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N422, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N424, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N426, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N428, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N430, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N432, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N434, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N436, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N438, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N440, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N442, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N444, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N446, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N448, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N450, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N452, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N454, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N456, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N458, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N460, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N462, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N464, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N466, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N468, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N470, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N472, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N411, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N413, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N415, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N417, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N419, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N421, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N423, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N425, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N427, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N429, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N431, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N433, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N435, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N437, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N439, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N441, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N443, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N445, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N447, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N449, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N451, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N453, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N455, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N457, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N459, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N461, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N463, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N465, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N467, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N469, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N471, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N473, 
         -- Connections to port 'Z'
         Z(0) => N481 );
   C12899_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_23_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_23_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_23_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_23_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_23_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_23_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_23_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_23_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_23_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_23_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_23_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_23_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_23_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_23_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_23_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_23_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_23_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_23_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_23_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_23_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_23_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_23_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_23_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_23_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_23_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_23_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_23_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_23_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_23_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_23_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_23_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_23_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_23_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_23_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_23_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_23_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_23_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_23_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_23_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_23_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_23_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_23_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_23_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_23_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_23_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_23_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_23_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_23_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_23_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_23_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_23_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_23_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_23_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_23_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_23_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_23_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_23_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_23_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_23_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_23_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_23_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_23_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_23_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_23_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N410, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N412, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N414, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N416, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N418, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N420, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N422, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N424, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N426, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N428, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N430, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N432, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N434, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N436, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N438, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N440, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N442, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N444, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N446, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N448, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N450, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N452, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N454, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N456, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N458, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N460, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N462, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N464, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N466, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N468, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N470, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N472, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N411, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N413, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N415, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N417, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N419, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N421, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N423, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N425, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N427, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N429, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N431, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N433, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N435, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N437, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N439, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N441, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N443, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N445, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N447, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N449, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N451, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N453, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N455, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N457, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N459, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N461, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N463, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N465, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N467, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N469, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N471, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N473, 
         -- Connections to port 'Z'
         Z(0) => N482 );
   C12900_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_22_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_22_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_22_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_22_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_22_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_22_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_22_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_22_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_22_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_22_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_22_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_22_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_22_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_22_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_22_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_22_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_22_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_22_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_22_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_22_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_22_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_22_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_22_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_22_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_22_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_22_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_22_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_22_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_22_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_22_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_22_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_22_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_22_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_22_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_22_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_22_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_22_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_22_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_22_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_22_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_22_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_22_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_22_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_22_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_22_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_22_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_22_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_22_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_22_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_22_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_22_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_22_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_22_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_22_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_22_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_22_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_22_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_22_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_22_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_22_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_22_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_22_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_22_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_22_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N410, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N412, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N414, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N416, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N418, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N420, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N422, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N424, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N426, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N428, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N430, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N432, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N434, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N436, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N438, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N440, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N442, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N444, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N446, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N448, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N450, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N452, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N454, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N456, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N458, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N460, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N462, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N464, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N466, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N468, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N470, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N472, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N411, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N413, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N415, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N417, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N419, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N421, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N423, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N425, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N427, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N429, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N431, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N433, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N435, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N437, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N439, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N441, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N443, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N445, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N447, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N449, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N451, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N453, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N455, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N457, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N459, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N461, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N463, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N465, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N467, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N469, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N471, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N473, 
         -- Connections to port 'Z'
         Z(0) => N483 );
   C12901_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_21_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_21_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_21_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_21_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_21_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_21_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_21_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_21_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_21_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_21_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_21_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_21_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_21_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_21_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_21_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_21_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_21_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_21_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_21_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_21_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_21_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_21_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_21_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_21_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_21_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_21_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_21_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_21_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_21_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_21_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_21_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_21_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_21_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_21_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_21_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_21_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_21_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_21_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_21_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_21_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_21_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_21_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_21_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_21_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_21_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_21_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_21_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_21_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_21_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_21_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_21_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_21_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_21_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_21_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_21_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_21_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_21_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_21_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_21_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_21_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_21_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_21_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_21_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_21_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N410, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N412, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N414, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N416, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N418, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N420, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N422, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N424, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N426, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N428, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N430, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N432, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N434, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N436, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N438, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N440, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N442, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N444, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N446, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N448, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N450, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N452, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N454, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N456, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N458, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N460, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N462, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N464, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N466, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N468, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N470, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N472, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N411, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N413, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N415, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N417, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N419, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N421, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N423, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N425, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N427, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N429, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N431, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N433, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N435, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N437, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N439, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N441, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N443, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N445, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N447, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N449, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N451, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N453, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N455, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N457, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N459, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N461, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N463, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N465, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N467, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N469, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N471, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N473, 
         -- Connections to port 'Z'
         Z(0) => N484 );
   C12902_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_20_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_20_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_20_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_20_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_20_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_20_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_20_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_20_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_20_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_20_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_20_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_20_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_20_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_20_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_20_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_20_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_20_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_20_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_20_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_20_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_20_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_20_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_20_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_20_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_20_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_20_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_20_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_20_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_20_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_20_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_20_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_20_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_20_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_20_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_20_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_20_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_20_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_20_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_20_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_20_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_20_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_20_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_20_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_20_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_20_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_20_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_20_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_20_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_20_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_20_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_20_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_20_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_20_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_20_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_20_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_20_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_20_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_20_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_20_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_20_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_20_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_20_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_20_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_20_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N410, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N412, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N414, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N416, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N418, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N420, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N422, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N424, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N426, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N428, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N430, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N432, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N434, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N436, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N438, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N440, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N442, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N444, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N446, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N448, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N450, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N452, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N454, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N456, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N458, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N460, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N462, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N464, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N466, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N468, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N470, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N472, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N411, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N413, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N415, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N417, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N419, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N421, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N423, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N425, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N427, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N429, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N431, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N433, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N435, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N437, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N439, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N441, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N443, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N445, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N447, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N449, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N451, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N453, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N455, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N457, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N459, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N461, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N463, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N465, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N467, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N469, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N471, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N473, 
         -- Connections to port 'Z'
         Z(0) => N485 );
   C12903_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_19_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_19_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_19_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_19_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_19_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_19_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_19_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_19_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_19_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_19_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_19_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_19_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_19_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_19_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_19_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_19_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_19_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_19_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_19_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_19_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_19_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_19_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_19_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_19_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_19_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_19_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_19_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_19_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_19_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_19_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_19_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_19_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_19_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_19_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_19_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_19_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_19_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_19_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_19_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_19_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_19_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_19_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_19_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_19_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_19_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_19_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_19_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_19_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_19_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_19_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_19_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_19_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_19_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_19_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_19_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_19_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_19_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_19_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_19_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_19_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_19_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_19_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_19_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_19_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N410, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N412, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N414, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N416, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N418, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N420, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N422, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N424, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N426, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N428, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N430, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N432, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N434, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N436, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N438, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N440, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N442, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N444, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N446, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N448, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N450, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N452, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N454, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N456, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N458, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N460, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N462, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N464, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N466, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N468, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N470, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N472, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N411, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N413, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N415, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N417, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N419, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N421, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N423, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N425, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N427, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N429, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N431, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N433, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N435, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N437, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N439, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N441, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N443, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N445, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N447, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N449, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N451, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N453, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N455, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N457, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N459, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N461, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N463, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N465, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N467, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N469, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N471, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N473, 
         -- Connections to port 'Z'
         Z(0) => N486 );
   C12904_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_18_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_18_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_18_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_18_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_18_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_18_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_18_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_18_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_18_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_18_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_18_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_18_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_18_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_18_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_18_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_18_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_18_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_18_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_18_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_18_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_18_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_18_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_18_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_18_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_18_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_18_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_18_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_18_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_18_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_18_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_18_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_18_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_18_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_18_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_18_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_18_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_18_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_18_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_18_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_18_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_18_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_18_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_18_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_18_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_18_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_18_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_18_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_18_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_18_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_18_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_18_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_18_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_18_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_18_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_18_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_18_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_18_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_18_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_18_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_18_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_18_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_18_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_18_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_18_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N410, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N412, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N414, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N416, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N418, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N420, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N422, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N424, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N426, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N428, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N430, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N432, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N434, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N436, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N438, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N440, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N442, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N444, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N446, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N448, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N450, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N452, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N454, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N456, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N458, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N460, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N462, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N464, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N466, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N468, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N470, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N472, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N411, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N413, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N415, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N417, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N419, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N421, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N423, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N425, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N427, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N429, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N431, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N433, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N435, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N437, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N439, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N441, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N443, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N445, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N447, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N449, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N451, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N453, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N455, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N457, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N459, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N461, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N463, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N465, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N467, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N469, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N471, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N473, 
         -- Connections to port 'Z'
         Z(0) => N487 );
   C12905_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_17_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_17_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_17_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_17_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_17_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_17_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_17_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_17_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_17_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_17_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_17_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_17_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_17_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_17_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_17_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_17_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_17_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_17_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_17_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_17_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_17_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_17_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_17_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_17_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_17_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_17_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_17_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_17_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_17_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_17_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_17_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_17_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_17_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_17_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_17_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_17_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_17_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_17_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_17_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_17_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_17_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_17_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_17_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_17_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_17_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_17_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_17_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_17_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_17_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_17_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_17_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_17_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_17_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_17_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_17_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_17_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_17_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_17_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_17_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_17_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_17_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_17_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_17_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_17_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N410, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N412, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N414, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N416, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N418, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N420, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N422, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N424, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N426, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N428, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N430, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N432, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N434, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N436, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N438, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N440, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N442, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N444, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N446, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N448, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N450, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N452, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N454, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N456, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N458, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N460, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N462, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N464, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N466, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N468, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N470, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N472, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N411, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N413, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N415, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N417, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N419, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N421, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N423, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N425, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N427, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N429, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N431, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N433, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N435, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N437, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N439, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N441, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N443, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N445, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N447, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N449, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N451, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N453, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N455, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N457, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N459, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N461, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N463, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N465, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N467, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N469, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N471, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N473, 
         -- Connections to port 'Z'
         Z(0) => N488 );
   C12906_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_16_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_16_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_16_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_16_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_16_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_16_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_16_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_16_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_16_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_16_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_16_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_16_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_16_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_16_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_16_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_16_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_16_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_16_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_16_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_16_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_16_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_16_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_16_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_16_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_16_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_16_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_16_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_16_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_16_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_16_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_16_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_16_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_16_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_16_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_16_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_16_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_16_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_16_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_16_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_16_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_16_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_16_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_16_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_16_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_16_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_16_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_16_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_16_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_16_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_16_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_16_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_16_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_16_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_16_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_16_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_16_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_16_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_16_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_16_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_16_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_16_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_16_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_16_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_16_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N410, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N412, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N414, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N416, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N418, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N420, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N422, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N424, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N426, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N428, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N430, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N432, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N434, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N436, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N438, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N440, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N442, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N444, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N446, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N448, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N450, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N452, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N454, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N456, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N458, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N460, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N462, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N464, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N466, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N468, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N470, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N472, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N411, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N413, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N415, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N417, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N419, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N421, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N423, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N425, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N427, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N429, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N431, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N433, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N435, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N437, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N439, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N441, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N443, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N445, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N447, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N449, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N451, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N453, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N455, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N457, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N459, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N461, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N463, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N465, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N467, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N469, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N471, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N473, 
         -- Connections to port 'Z'
         Z(0) => N489 );
   C12907_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_15_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_15_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_15_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_15_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_15_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_15_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_15_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_15_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_15_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_15_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_15_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_15_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_15_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_15_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_15_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_15_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_15_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_15_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_15_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_15_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_15_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_15_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_15_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_15_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_15_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_15_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_15_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_15_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_15_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_15_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_15_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_15_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_15_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_15_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_15_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_15_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_15_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_15_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_15_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_15_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_15_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_15_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_15_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_15_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_15_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_15_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_15_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_15_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_15_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_15_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_15_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_15_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_15_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_15_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_15_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_15_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_15_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_15_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_15_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_15_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_15_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_15_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_15_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_15_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N410, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N412, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N414, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N416, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N418, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N420, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N422, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N424, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N426, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N428, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N430, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N432, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N434, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N436, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N438, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N440, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N442, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N444, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N446, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N448, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N450, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N452, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N454, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N456, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N458, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N460, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N462, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N464, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N466, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N468, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N470, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N472, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N411, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N413, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N415, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N417, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N419, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N421, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N423, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N425, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N427, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N429, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N431, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N433, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N435, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N437, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N439, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N441, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N443, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N445, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N447, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N449, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N451, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N453, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N455, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N457, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N459, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N461, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N463, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N465, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N467, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N469, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N471, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N473, 
         -- Connections to port 'Z'
         Z(0) => N490 );
   C12908_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_14_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_14_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_14_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_14_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_14_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_14_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_14_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_14_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_14_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_14_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_14_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_14_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_14_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_14_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_14_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_14_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_14_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_14_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_14_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_14_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_14_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_14_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_14_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_14_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_14_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_14_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_14_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_14_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_14_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_14_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_14_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_14_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_14_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_14_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_14_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_14_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_14_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_14_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_14_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_14_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_14_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_14_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_14_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_14_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_14_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_14_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_14_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_14_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_14_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_14_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_14_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_14_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_14_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_14_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_14_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_14_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_14_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_14_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_14_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_14_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_14_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_14_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_14_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_14_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N410, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N412, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N414, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N416, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N418, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N420, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N422, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N424, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N426, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N428, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N430, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N432, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N434, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N436, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N438, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N440, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N442, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N444, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N446, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N448, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N450, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N452, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N454, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N456, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N458, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N460, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N462, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N464, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N466, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N468, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N470, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N472, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N411, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N413, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N415, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N417, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N419, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N421, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N423, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N425, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N427, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N429, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N431, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N433, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N435, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N437, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N439, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N441, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N443, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N445, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N447, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N449, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N451, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N453, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N455, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N457, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N459, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N461, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N463, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N465, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N467, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N469, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N471, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N473, 
         -- Connections to port 'Z'
         Z(0) => N491 );
   C12909_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_13_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_13_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_13_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_13_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_13_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_13_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_13_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_13_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_13_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_13_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_13_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_13_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_13_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_13_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_13_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_13_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_13_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_13_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_13_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_13_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_13_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_13_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_13_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_13_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_13_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_13_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_13_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_13_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_13_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_13_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_13_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_13_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_13_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_13_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_13_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_13_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_13_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_13_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_13_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_13_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_13_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_13_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_13_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_13_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_13_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_13_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_13_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_13_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_13_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_13_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_13_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_13_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_13_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_13_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_13_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_13_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_13_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_13_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_13_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_13_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_13_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_13_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_13_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_13_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N410, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N412, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N414, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N416, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N418, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N420, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N422, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N424, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N426, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N428, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N430, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N432, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N434, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N436, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N438, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N440, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N442, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N444, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N446, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N448, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N450, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N452, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N454, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N456, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N458, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N460, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N462, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N464, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N466, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N468, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N470, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N472, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N411, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N413, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N415, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N417, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N419, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N421, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N423, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N425, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N427, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N429, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N431, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N433, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N435, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N437, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N439, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N441, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N443, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N445, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N447, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N449, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N451, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N453, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N455, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N457, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N459, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N461, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N463, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N465, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N467, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N469, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N471, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N473, 
         -- Connections to port 'Z'
         Z(0) => N492 );
   C12910_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_12_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_12_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_12_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_12_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_12_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_12_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_12_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_12_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_12_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_12_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_12_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_12_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_12_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_12_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_12_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_12_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_12_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_12_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_12_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_12_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_12_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_12_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_12_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_12_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_12_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_12_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_12_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_12_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_12_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_12_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_12_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_12_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_12_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_12_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_12_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_12_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_12_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_12_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_12_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_12_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_12_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_12_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_12_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_12_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_12_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_12_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_12_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_12_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_12_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_12_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_12_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_12_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_12_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_12_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_12_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_12_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_12_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_12_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_12_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_12_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_12_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_12_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_12_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_12_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N410, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N412, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N414, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N416, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N418, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N420, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N422, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N424, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N426, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N428, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N430, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N432, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N434, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N436, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N438, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N440, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N442, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N444, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N446, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N448, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N450, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N452, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N454, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N456, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N458, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N460, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N462, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N464, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N466, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N468, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N470, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N472, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N411, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N413, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N415, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N417, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N419, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N421, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N423, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N425, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N427, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N429, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N431, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N433, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N435, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N437, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N439, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N441, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N443, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N445, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N447, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N449, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N451, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N453, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N455, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N457, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N459, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N461, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N463, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N465, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N467, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N469, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N471, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N473, 
         -- Connections to port 'Z'
         Z(0) => N493 );
   C12911_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_11_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_11_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_11_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_11_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_11_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_11_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_11_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_11_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_11_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_11_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_11_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_11_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_11_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_11_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_11_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_11_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_11_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_11_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_11_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_11_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_11_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_11_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_11_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_11_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_11_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_11_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_11_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_11_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_11_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_11_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_11_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_11_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_11_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_11_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_11_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_11_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_11_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_11_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_11_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_11_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_11_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_11_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_11_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_11_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_11_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_11_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_11_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_11_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_11_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_11_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_11_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_11_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_11_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_11_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_11_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_11_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_11_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_11_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_11_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_11_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_11_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_11_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_11_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_11_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N410, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N412, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N414, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N416, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N418, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N420, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N422, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N424, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N426, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N428, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N430, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N432, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N434, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N436, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N438, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N440, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N442, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N444, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N446, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N448, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N450, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N452, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N454, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N456, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N458, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N460, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N462, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N464, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N466, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N468, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N470, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N472, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N411, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N413, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N415, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N417, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N419, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N421, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N423, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N425, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N427, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N429, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N431, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N433, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N435, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N437, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N439, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N441, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N443, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N445, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N447, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N449, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N451, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N453, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N455, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N457, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N459, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N461, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N463, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N465, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N467, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N469, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N471, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N473, 
         -- Connections to port 'Z'
         Z(0) => N494 );
   C12912_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_10_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_10_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_10_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_10_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_10_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_10_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_10_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_10_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_10_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_10_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_10_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_10_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_10_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_10_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_10_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_10_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_10_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_10_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_10_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_10_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_10_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_10_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_10_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_10_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_10_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_10_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_10_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_10_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_10_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_10_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_10_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_10_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_10_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_10_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_10_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_10_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_10_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_10_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_10_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_10_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_10_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_10_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_10_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_10_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_10_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_10_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_10_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_10_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_10_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_10_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_10_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_10_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_10_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_10_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_10_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_10_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_10_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_10_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_10_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_10_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_10_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_10_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_10_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_10_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N410, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N412, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N414, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N416, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N418, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N420, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N422, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N424, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N426, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N428, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N430, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N432, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N434, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N436, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N438, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N440, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N442, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N444, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N446, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N448, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N450, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N452, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N454, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N456, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N458, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N460, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N462, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N464, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N466, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N468, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N470, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N472, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N411, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N413, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N415, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N417, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N419, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N421, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N423, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N425, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N427, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N429, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N431, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N433, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N435, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N437, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N439, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N441, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N443, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N445, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N447, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N449, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N451, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N453, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N455, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N457, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N459, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N461, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N463, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N465, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N467, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N469, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N471, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N473, 
         -- Connections to port 'Z'
         Z(0) => N495 );
   C12913_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_9_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_9_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_9_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_9_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_9_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_9_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_9_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_9_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_9_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_9_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_9_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_9_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_9_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_9_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_9_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_9_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_9_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_9_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_9_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_9_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_9_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_9_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_9_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_9_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_9_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_9_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_9_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_9_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_9_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_9_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_9_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_9_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_9_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_9_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_9_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_9_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_9_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_9_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_9_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_9_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_9_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_9_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_9_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_9_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_9_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_9_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_9_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_9_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_9_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_9_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_9_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_9_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_9_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_9_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_9_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_9_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_9_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_9_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_9_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_9_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_9_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_9_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_9_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_9_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N410, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N412, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N414, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N416, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N418, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N420, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N422, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N424, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N426, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N428, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N430, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N432, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N434, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N436, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N438, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N440, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N442, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N444, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N446, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N448, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N450, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N452, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N454, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N456, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N458, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N460, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N462, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N464, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N466, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N468, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N470, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N472, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N411, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N413, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N415, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N417, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N419, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N421, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N423, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N425, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N427, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N429, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N431, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N433, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N435, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N437, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N439, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N441, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N443, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N445, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N447, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N449, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N451, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N453, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N455, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N457, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N459, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N461, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N463, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N465, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N467, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N469, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N471, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N473, 
         -- Connections to port 'Z'
         Z(0) => N496 );
   C12914_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_8_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_8_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_8_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_8_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_8_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_8_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_8_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_8_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_8_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_8_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_8_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_8_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_8_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_8_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_8_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_8_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_8_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_8_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_8_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_8_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_8_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_8_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_8_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_8_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_8_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_8_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_8_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_8_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_8_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_8_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_8_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_8_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_8_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_8_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_8_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_8_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_8_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_8_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_8_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_8_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_8_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_8_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_8_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_8_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_8_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_8_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_8_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_8_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_8_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_8_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_8_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_8_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_8_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_8_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_8_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_8_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_8_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_8_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_8_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_8_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_8_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_8_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_8_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_8_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N410, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N412, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N414, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N416, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N418, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N420, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N422, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N424, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N426, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N428, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N430, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N432, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N434, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N436, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N438, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N440, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N442, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N444, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N446, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N448, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N450, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N452, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N454, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N456, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N458, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N460, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N462, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N464, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N466, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N468, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N470, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N472, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N411, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N413, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N415, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N417, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N419, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N421, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N423, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N425, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N427, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N429, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N431, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N433, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N435, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N437, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N439, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N441, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N443, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N445, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N447, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N449, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N451, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N453, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N455, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N457, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N459, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N461, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N463, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N465, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N467, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N469, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N471, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N473, 
         -- Connections to port 'Z'
         Z(0) => N497 );
   C12915_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_7_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_7_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_7_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_7_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_7_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_7_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_7_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_7_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_7_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_7_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_7_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_7_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_7_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_7_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_7_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_7_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_7_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_7_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_7_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_7_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_7_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_7_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_7_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_7_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_7_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_7_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_7_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_7_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_7_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_7_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_7_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_7_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_7_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_7_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_7_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_7_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_7_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_7_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_7_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_7_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_7_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_7_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_7_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_7_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_7_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_7_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_7_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_7_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_7_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_7_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_7_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_7_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_7_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_7_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_7_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_7_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_7_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_7_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_7_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_7_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_7_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_7_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_7_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_7_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N410, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N412, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N414, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N416, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N418, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N420, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N422, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N424, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N426, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N428, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N430, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N432, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N434, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N436, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N438, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N440, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N442, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N444, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N446, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N448, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N450, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N452, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N454, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N456, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N458, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N460, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N462, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N464, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N466, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N468, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N470, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N472, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N411, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N413, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N415, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N417, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N419, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N421, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N423, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N425, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N427, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N429, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N431, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N433, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N435, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N437, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N439, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N441, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N443, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N445, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N447, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N449, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N451, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N453, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N455, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N457, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N459, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N461, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N463, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N465, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N467, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N469, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N471, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N473, 
         -- Connections to port 'Z'
         Z(0) => N498 );
   C12916_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_6_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_6_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_6_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_6_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_6_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_6_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_6_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_6_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_6_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_6_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_6_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_6_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_6_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_6_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_6_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_6_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_6_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_6_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_6_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_6_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_6_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_6_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_6_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_6_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_6_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_6_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_6_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_6_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_6_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_6_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_6_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_6_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_6_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_6_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_6_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_6_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_6_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_6_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_6_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_6_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_6_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_6_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_6_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_6_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_6_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_6_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_6_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_6_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_6_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_6_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_6_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_6_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_6_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_6_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_6_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_6_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_6_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_6_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_6_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_6_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_6_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_6_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_6_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_6_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N410, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N412, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N414, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N416, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N418, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N420, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N422, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N424, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N426, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N428, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N430, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N432, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N434, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N436, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N438, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N440, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N442, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N444, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N446, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N448, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N450, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N452, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N454, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N456, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N458, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N460, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N462, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N464, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N466, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N468, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N470, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N472, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N411, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N413, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N415, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N417, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N419, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N421, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N423, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N425, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N427, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N429, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N431, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N433, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N435, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N437, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N439, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N441, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N443, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N445, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N447, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N449, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N451, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N453, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N455, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N457, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N459, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N461, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N463, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N465, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N467, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N469, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N471, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N473, 
         -- Connections to port 'Z'
         Z(0) => N499 );
   C12917_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_5_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_5_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_5_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_5_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_5_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_5_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_5_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_5_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_5_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_5_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_5_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_5_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_5_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_5_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_5_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_5_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_5_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_5_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_5_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_5_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_5_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_5_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_5_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_5_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_5_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_5_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_5_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_5_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_5_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_5_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_5_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_5_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_5_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_5_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_5_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_5_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_5_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_5_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_5_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_5_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_5_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_5_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_5_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_5_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_5_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_5_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_5_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_5_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_5_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_5_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_5_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_5_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_5_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_5_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_5_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_5_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_5_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_5_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_5_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_5_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_5_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_5_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_5_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_5_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N410, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N412, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N414, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N416, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N418, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N420, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N422, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N424, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N426, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N428, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N430, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N432, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N434, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N436, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N438, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N440, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N442, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N444, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N446, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N448, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N450, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N452, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N454, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N456, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N458, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N460, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N462, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N464, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N466, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N468, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N470, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N472, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N411, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N413, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N415, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N417, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N419, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N421, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N423, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N425, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N427, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N429, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N431, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N433, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N435, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N437, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N439, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N441, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N443, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N445, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N447, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N449, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N451, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N453, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N455, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N457, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N459, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N461, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N463, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N465, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N467, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N469, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N471, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N473, 
         -- Connections to port 'Z'
         Z(0) => N500 );
   C12918_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_4_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_4_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_4_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_4_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_4_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_4_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_4_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_4_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_4_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_4_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_4_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_4_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_4_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_4_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_4_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_4_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_4_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_4_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_4_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_4_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_4_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_4_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_4_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_4_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_4_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_4_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_4_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_4_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_4_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_4_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_4_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_4_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_4_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_4_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_4_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_4_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_4_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_4_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_4_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_4_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_4_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_4_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_4_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_4_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_4_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_4_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_4_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_4_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_4_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_4_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_4_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_4_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_4_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_4_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_4_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_4_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_4_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_4_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_4_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_4_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_4_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_4_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_4_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_4_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N410, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N412, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N414, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N416, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N418, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N420, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N422, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N424, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N426, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N428, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N430, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N432, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N434, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N436, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N438, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N440, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N442, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N444, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N446, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N448, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N450, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N452, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N454, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N456, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N458, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N460, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N462, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N464, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N466, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N468, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N470, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N472, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N411, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N413, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N415, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N417, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N419, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N421, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N423, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N425, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N427, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N429, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N431, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N433, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N435, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N437, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N439, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N441, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N443, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N445, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N447, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N449, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N451, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N453, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N455, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N457, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N459, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N461, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N463, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N465, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N467, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N469, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N471, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N473, 
         -- Connections to port 'Z'
         Z(0) => N501 );
   C12919_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_3_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_3_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_3_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_3_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_3_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_3_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_3_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_3_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_3_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_3_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_3_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_3_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_3_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_3_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_3_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_3_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_3_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_3_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_3_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_3_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_3_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_3_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_3_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_3_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_3_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_3_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_3_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_3_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_3_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_3_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_3_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_3_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_3_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_3_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_3_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_3_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_3_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_3_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_3_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_3_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_3_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_3_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_3_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_3_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_3_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_3_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_3_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_3_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_3_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_3_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_3_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_3_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_3_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_3_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_3_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_3_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_3_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_3_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_3_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_3_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_3_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_3_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_3_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_3_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N410, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N412, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N414, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N416, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N418, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N420, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N422, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N424, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N426, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N428, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N430, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N432, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N434, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N436, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N438, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N440, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N442, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N444, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N446, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N448, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N450, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N452, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N454, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N456, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N458, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N460, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N462, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N464, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N466, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N468, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N470, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N472, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N411, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N413, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N415, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N417, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N419, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N421, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N423, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N425, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N427, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N429, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N431, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N433, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N435, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N437, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N439, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N441, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N443, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N445, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N447, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N449, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N451, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N453, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N455, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N457, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N459, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N461, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N463, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N465, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N467, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N469, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N471, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N473, 
         -- Connections to port 'Z'
         Z(0) => N502 );
   C12920_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_2_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_2_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_2_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_2_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_2_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_2_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_2_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_2_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_2_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_2_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_2_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_2_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_2_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_2_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_2_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_2_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_2_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_2_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_2_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_2_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_2_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_2_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_2_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_2_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_2_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_2_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_2_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_2_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_2_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_2_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_2_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_2_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_2_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_2_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_2_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_2_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_2_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_2_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_2_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_2_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_2_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_2_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_2_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_2_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_2_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_2_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_2_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_2_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_2_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_2_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_2_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_2_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_2_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_2_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_2_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_2_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_2_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_2_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_2_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_2_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_2_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_2_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_2_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_2_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N410, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N412, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N414, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N416, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N418, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N420, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N422, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N424, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N426, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N428, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N430, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N432, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N434, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N436, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N438, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N440, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N442, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N444, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N446, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N448, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N450, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N452, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N454, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N456, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N458, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N460, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N462, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N464, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N466, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N468, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N470, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N472, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N411, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N413, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N415, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N417, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N419, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N421, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N423, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N425, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N427, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N429, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N431, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N433, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N435, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N437, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N439, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N441, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N443, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N445, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N447, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N449, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N451, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N453, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N455, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N457, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N459, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N461, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N463, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N465, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N467, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N469, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N471, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N473, 
         -- Connections to port 'Z'
         Z(0) => N503 );
   C12921_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_1_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_1_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_1_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_1_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_1_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_1_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_1_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_1_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_1_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_1_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_1_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_1_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_1_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_1_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_1_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_1_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_1_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_1_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_1_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_1_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_1_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_1_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_1_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_1_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_1_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_1_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_1_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_1_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_1_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_1_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_1_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_1_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_1_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_1_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_1_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_1_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_1_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_1_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_1_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_1_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_1_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_1_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_1_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_1_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_1_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_1_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_1_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_1_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_1_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_1_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_1_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_1_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_1_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_1_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_1_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_1_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_1_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_1_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_1_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_1_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_1_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_1_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_1_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_1_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N410, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N412, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N414, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N416, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N418, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N420, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N422, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N424, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N426, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N428, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N430, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N432, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N434, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N436, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N438, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N440, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N442, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N444, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N446, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N448, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N450, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N452, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N454, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N456, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N458, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N460, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N462, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N464, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N466, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N468, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N470, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N472, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N411, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N413, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N415, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N417, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N419, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N421, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N423, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N425, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N427, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N429, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N431, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N433, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N435, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N437, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N439, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N441, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N443, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N445, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N447, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N449, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N451, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N453, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N455, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N457, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N459, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N461, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N463, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N465, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N467, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N469, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N471, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N473, 
         -- Connections to port 'Z'
         Z(0) => N504 );
   C12922_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_0_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_0_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_0_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_0_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_0_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_0_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_0_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_0_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_0_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_0_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_0_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_0_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_0_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_0_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_0_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_0_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_0_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_0_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_0_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_0_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_0_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_0_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_0_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_0_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_0_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_0_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_0_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_0_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_0_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_0_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_0_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_0_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_0_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_0_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_0_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_0_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_0_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_0_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_0_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_0_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_0_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_0_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_0_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_0_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_0_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_0_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_0_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_0_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_0_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_0_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_0_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_0_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_0_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_0_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_0_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_0_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_0_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_0_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_0_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_0_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_0_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_0_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N410, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N412, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N414, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N416, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N418, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N420, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N422, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N424, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N426, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N428, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N430, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N432, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N434, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N436, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N438, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N440, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N442, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N444, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N446, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N448, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N450, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N452, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N454, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N456, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N458, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N460, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N462, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N464, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N466, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N468, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N470, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N472, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N411, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N413, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N415, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N417, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N419, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N421, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N423, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N425, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N427, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N429, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N431, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N433, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N435, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N437, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N439, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N441, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N443, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N445, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N447, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N449, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N451, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N453, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N455, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N457, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N459, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N461, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N463, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N465, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N467, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N469, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N471, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N473, 
         -- Connections to port 'Z'
         Z(0) => N505 );
   C13059_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_31_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_31_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_31_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_31_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_31_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_31_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_31_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_31_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_31_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_31_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_31_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_31_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_31_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_31_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_31_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_31_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_31_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_31_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_31_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_31_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_31_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_31_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_31_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_31_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_31_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_31_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_31_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_31_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_31_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_31_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_31_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_31_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_31_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_31_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_31_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_31_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_31_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_31_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_31_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_31_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_31_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_31_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_31_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_31_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_31_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_31_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_31_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_31_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_31_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_31_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_31_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_31_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_31_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_31_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_31_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_31_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_31_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_31_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_31_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_31_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_31_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_31_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_31_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_31_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N248, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N252, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N254, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N256, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N258, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N260, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N262, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N264, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N266, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N268, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N270, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N272, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N274, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N276, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N278, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N280, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N282, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N284, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N286, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N288, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N290, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N292, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N294, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N296, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N298, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N300, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N302, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N304, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N306, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N308, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N310, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N249, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N251, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N253, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N255, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N257, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N259, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N261, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N263, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N265, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N267, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N269, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N271, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N273, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N275, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N277, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N279, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N281, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N283, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N285, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N287, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N289, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N291, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N293, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N295, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N297, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N299, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N301, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N303, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N305, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N307, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N309, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N311, 
         -- Connections to port 'Z'
         Z(0) => N507 );
   C13060_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_30_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_30_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_30_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_30_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_30_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_30_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_30_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_30_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_30_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_30_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_30_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_30_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_30_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_30_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_30_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_30_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_30_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_30_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_30_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_30_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_30_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_30_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_30_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_30_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_30_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_30_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_30_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_30_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_30_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_30_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_30_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_30_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_30_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_30_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_30_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_30_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_30_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_30_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_30_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_30_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_30_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_30_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_30_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_30_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_30_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_30_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_30_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_30_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_30_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_30_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_30_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_30_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_30_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_30_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_30_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_30_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_30_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_30_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_30_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_30_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_30_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_30_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_30_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_30_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N248, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N252, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N254, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N256, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N258, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N260, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N262, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N264, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N266, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N268, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N270, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N272, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N274, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N276, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N278, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N280, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N282, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N284, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N286, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N288, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N290, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N292, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N294, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N296, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N298, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N300, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N302, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N304, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N306, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N308, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N310, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N249, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N251, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N253, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N255, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N257, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N259, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N261, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N263, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N265, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N267, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N269, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N271, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N273, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N275, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N277, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N279, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N281, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N283, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N285, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N287, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N289, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N291, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N293, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N295, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N297, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N299, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N301, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N303, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N305, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N307, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N309, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N311, 
         -- Connections to port 'Z'
         Z(0) => N508 );
   C13061_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_29_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_29_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_29_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_29_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_29_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_29_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_29_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_29_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_29_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_29_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_29_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_29_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_29_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_29_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_29_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_29_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_29_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_29_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_29_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_29_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_29_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_29_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_29_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_29_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_29_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_29_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_29_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_29_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_29_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_29_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_29_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_29_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_29_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_29_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_29_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_29_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_29_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_29_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_29_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_29_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_29_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_29_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_29_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_29_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_29_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_29_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_29_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_29_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_29_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_29_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_29_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_29_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_29_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_29_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_29_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_29_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_29_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_29_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_29_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_29_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_29_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_29_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_29_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_29_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N248, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N252, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N254, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N256, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N258, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N260, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N262, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N264, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N266, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N268, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N270, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N272, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N274, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N276, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N278, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N280, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N282, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N284, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N286, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N288, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N290, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N292, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N294, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N296, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N298, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N300, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N302, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N304, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N306, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N308, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N310, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N249, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N251, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N253, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N255, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N257, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N259, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N261, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N263, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N265, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N267, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N269, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N271, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N273, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N275, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N277, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N279, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N281, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N283, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N285, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N287, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N289, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N291, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N293, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N295, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N297, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N299, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N301, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N303, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N305, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N307, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N309, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N311, 
         -- Connections to port 'Z'
         Z(0) => N509 );
   C13062_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_28_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_28_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_28_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_28_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_28_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_28_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_28_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_28_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_28_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_28_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_28_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_28_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_28_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_28_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_28_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_28_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_28_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_28_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_28_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_28_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_28_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_28_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_28_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_28_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_28_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_28_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_28_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_28_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_28_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_28_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_28_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_28_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_28_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_28_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_28_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_28_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_28_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_28_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_28_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_28_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_28_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_28_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_28_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_28_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_28_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_28_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_28_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_28_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_28_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_28_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_28_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_28_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_28_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_28_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_28_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_28_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_28_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_28_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_28_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_28_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_28_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_28_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_28_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_28_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N248, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N252, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N254, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N256, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N258, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N260, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N262, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N264, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N266, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N268, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N270, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N272, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N274, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N276, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N278, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N280, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N282, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N284, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N286, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N288, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N290, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N292, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N294, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N296, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N298, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N300, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N302, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N304, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N306, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N308, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N310, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N249, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N251, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N253, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N255, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N257, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N259, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N261, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N263, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N265, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N267, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N269, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N271, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N273, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N275, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N277, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N279, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N281, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N283, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N285, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N287, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N289, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N291, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N293, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N295, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N297, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N299, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N301, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N303, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N305, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N307, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N309, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N311, 
         -- Connections to port 'Z'
         Z(0) => N510 );
   C13063_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_27_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_27_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_27_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_27_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_27_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_27_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_27_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_27_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_27_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_27_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_27_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_27_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_27_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_27_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_27_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_27_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_27_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_27_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_27_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_27_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_27_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_27_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_27_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_27_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_27_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_27_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_27_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_27_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_27_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_27_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_27_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_27_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_27_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_27_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_27_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_27_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_27_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_27_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_27_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_27_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_27_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_27_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_27_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_27_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_27_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_27_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_27_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_27_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_27_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_27_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_27_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_27_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_27_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_27_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_27_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_27_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_27_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_27_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_27_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_27_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_27_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_27_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_27_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_27_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N248, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N252, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N254, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N256, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N258, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N260, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N262, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N264, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N266, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N268, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N270, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N272, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N274, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N276, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N278, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N280, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N282, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N284, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N286, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N288, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N290, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N292, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N294, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N296, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N298, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N300, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N302, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N304, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N306, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N308, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N310, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N249, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N251, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N253, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N255, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N257, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N259, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N261, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N263, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N265, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N267, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N269, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N271, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N273, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N275, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N277, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N279, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N281, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N283, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N285, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N287, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N289, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N291, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N293, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N295, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N297, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N299, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N301, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N303, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N305, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N307, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N309, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N311, 
         -- Connections to port 'Z'
         Z(0) => N511 );
   C13064_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_26_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_26_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_26_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_26_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_26_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_26_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_26_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_26_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_26_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_26_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_26_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_26_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_26_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_26_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_26_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_26_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_26_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_26_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_26_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_26_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_26_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_26_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_26_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_26_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_26_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_26_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_26_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_26_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_26_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_26_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_26_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_26_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_26_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_26_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_26_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_26_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_26_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_26_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_26_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_26_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_26_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_26_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_26_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_26_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_26_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_26_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_26_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_26_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_26_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_26_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_26_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_26_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_26_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_26_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_26_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_26_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_26_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_26_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_26_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_26_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_26_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_26_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_26_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_26_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N248, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N252, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N254, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N256, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N258, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N260, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N262, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N264, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N266, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N268, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N270, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N272, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N274, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N276, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N278, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N280, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N282, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N284, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N286, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N288, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N290, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N292, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N294, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N296, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N298, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N300, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N302, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N304, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N306, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N308, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N310, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N249, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N251, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N253, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N255, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N257, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N259, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N261, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N263, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N265, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N267, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N269, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N271, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N273, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N275, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N277, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N279, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N281, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N283, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N285, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N287, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N289, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N291, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N293, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N295, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N297, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N299, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N301, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N303, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N305, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N307, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N309, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N311, 
         -- Connections to port 'Z'
         Z(0) => N512 );
   C13065_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_25_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_25_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_25_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_25_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_25_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_25_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_25_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_25_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_25_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_25_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_25_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_25_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_25_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_25_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_25_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_25_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_25_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_25_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_25_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_25_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_25_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_25_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_25_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_25_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_25_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_25_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_25_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_25_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_25_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_25_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_25_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_25_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_25_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_25_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_25_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_25_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_25_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_25_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_25_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_25_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_25_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_25_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_25_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_25_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_25_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_25_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_25_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_25_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_25_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_25_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_25_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_25_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_25_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_25_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_25_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_25_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_25_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_25_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_25_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_25_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_25_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_25_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_25_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_25_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N248, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N252, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N254, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N256, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N258, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N260, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N262, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N264, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N266, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N268, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N270, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N272, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N274, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N276, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N278, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N280, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N282, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N284, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N286, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N288, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N290, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N292, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N294, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N296, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N298, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N300, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N302, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N304, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N306, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N308, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N310, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N249, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N251, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N253, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N255, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N257, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N259, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N261, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N263, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N265, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N267, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N269, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N271, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N273, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N275, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N277, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N279, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N281, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N283, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N285, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N287, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N289, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N291, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N293, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N295, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N297, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N299, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N301, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N303, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N305, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N307, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N309, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N311, 
         -- Connections to port 'Z'
         Z(0) => N513 );
   C13066_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_24_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_24_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_24_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_24_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_24_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_24_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_24_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_24_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_24_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_24_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_24_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_24_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_24_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_24_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_24_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_24_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_24_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_24_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_24_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_24_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_24_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_24_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_24_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_24_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_24_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_24_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_24_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_24_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_24_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_24_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_24_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_24_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_24_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_24_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_24_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_24_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_24_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_24_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_24_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_24_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_24_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_24_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_24_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_24_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_24_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_24_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_24_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_24_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_24_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_24_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_24_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_24_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_24_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_24_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_24_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_24_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_24_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_24_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_24_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_24_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_24_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_24_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_24_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_24_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N248, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N252, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N254, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N256, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N258, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N260, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N262, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N264, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N266, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N268, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N270, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N272, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N274, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N276, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N278, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N280, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N282, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N284, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N286, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N288, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N290, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N292, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N294, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N296, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N298, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N300, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N302, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N304, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N306, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N308, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N310, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N249, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N251, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N253, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N255, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N257, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N259, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N261, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N263, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N265, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N267, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N269, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N271, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N273, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N275, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N277, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N279, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N281, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N283, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N285, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N287, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N289, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N291, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N293, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N295, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N297, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N299, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N301, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N303, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N305, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N307, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N309, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N311, 
         -- Connections to port 'Z'
         Z(0) => N514 );
   C13067_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_23_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_23_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_23_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_23_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_23_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_23_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_23_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_23_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_23_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_23_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_23_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_23_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_23_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_23_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_23_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_23_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_23_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_23_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_23_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_23_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_23_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_23_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_23_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_23_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_23_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_23_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_23_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_23_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_23_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_23_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_23_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_23_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_23_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_23_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_23_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_23_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_23_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_23_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_23_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_23_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_23_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_23_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_23_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_23_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_23_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_23_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_23_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_23_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_23_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_23_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_23_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_23_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_23_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_23_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_23_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_23_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_23_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_23_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_23_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_23_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_23_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_23_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_23_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_23_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N248, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N252, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N254, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N256, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N258, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N260, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N262, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N264, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N266, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N268, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N270, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N272, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N274, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N276, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N278, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N280, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N282, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N284, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N286, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N288, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N290, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N292, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N294, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N296, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N298, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N300, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N302, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N304, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N306, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N308, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N310, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N249, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N251, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N253, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N255, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N257, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N259, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N261, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N263, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N265, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N267, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N269, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N271, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N273, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N275, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N277, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N279, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N281, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N283, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N285, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N287, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N289, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N291, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N293, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N295, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N297, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N299, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N301, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N303, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N305, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N307, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N309, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N311, 
         -- Connections to port 'Z'
         Z(0) => N515 );
   C13068_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_22_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_22_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_22_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_22_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_22_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_22_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_22_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_22_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_22_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_22_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_22_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_22_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_22_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_22_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_22_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_22_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_22_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_22_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_22_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_22_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_22_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_22_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_22_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_22_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_22_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_22_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_22_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_22_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_22_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_22_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_22_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_22_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_22_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_22_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_22_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_22_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_22_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_22_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_22_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_22_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_22_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_22_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_22_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_22_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_22_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_22_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_22_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_22_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_22_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_22_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_22_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_22_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_22_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_22_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_22_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_22_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_22_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_22_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_22_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_22_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_22_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_22_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_22_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_22_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N248, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N252, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N254, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N256, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N258, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N260, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N262, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N264, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N266, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N268, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N270, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N272, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N274, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N276, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N278, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N280, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N282, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N284, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N286, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N288, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N290, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N292, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N294, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N296, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N298, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N300, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N302, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N304, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N306, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N308, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N310, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N249, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N251, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N253, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N255, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N257, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N259, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N261, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N263, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N265, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N267, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N269, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N271, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N273, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N275, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N277, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N279, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N281, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N283, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N285, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N287, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N289, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N291, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N293, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N295, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N297, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N299, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N301, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N303, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N305, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N307, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N309, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N311, 
         -- Connections to port 'Z'
         Z(0) => N516 );
   C13069_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_21_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_21_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_21_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_21_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_21_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_21_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_21_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_21_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_21_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_21_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_21_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_21_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_21_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_21_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_21_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_21_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_21_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_21_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_21_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_21_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_21_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_21_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_21_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_21_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_21_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_21_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_21_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_21_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_21_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_21_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_21_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_21_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_21_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_21_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_21_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_21_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_21_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_21_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_21_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_21_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_21_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_21_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_21_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_21_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_21_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_21_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_21_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_21_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_21_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_21_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_21_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_21_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_21_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_21_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_21_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_21_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_21_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_21_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_21_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_21_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_21_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_21_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_21_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_21_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N248, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N252, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N254, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N256, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N258, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N260, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N262, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N264, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N266, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N268, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N270, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N272, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N274, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N276, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N278, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N280, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N282, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N284, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N286, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N288, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N290, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N292, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N294, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N296, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N298, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N300, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N302, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N304, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N306, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N308, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N310, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N249, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N251, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N253, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N255, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N257, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N259, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N261, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N263, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N265, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N267, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N269, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N271, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N273, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N275, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N277, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N279, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N281, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N283, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N285, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N287, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N289, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N291, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N293, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N295, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N297, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N299, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N301, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N303, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N305, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N307, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N309, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N311, 
         -- Connections to port 'Z'
         Z(0) => N517 );
   C13070_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_20_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_20_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_20_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_20_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_20_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_20_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_20_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_20_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_20_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_20_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_20_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_20_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_20_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_20_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_20_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_20_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_20_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_20_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_20_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_20_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_20_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_20_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_20_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_20_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_20_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_20_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_20_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_20_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_20_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_20_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_20_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_20_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_20_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_20_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_20_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_20_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_20_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_20_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_20_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_20_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_20_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_20_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_20_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_20_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_20_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_20_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_20_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_20_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_20_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_20_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_20_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_20_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_20_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_20_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_20_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_20_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_20_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_20_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_20_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_20_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_20_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_20_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_20_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_20_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N248, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N252, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N254, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N256, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N258, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N260, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N262, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N264, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N266, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N268, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N270, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N272, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N274, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N276, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N278, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N280, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N282, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N284, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N286, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N288, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N290, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N292, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N294, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N296, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N298, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N300, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N302, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N304, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N306, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N308, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N310, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N249, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N251, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N253, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N255, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N257, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N259, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N261, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N263, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N265, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N267, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N269, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N271, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N273, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N275, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N277, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N279, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N281, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N283, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N285, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N287, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N289, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N291, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N293, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N295, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N297, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N299, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N301, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N303, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N305, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N307, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N309, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N311, 
         -- Connections to port 'Z'
         Z(0) => N518 );
   C13071_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_19_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_19_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_19_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_19_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_19_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_19_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_19_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_19_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_19_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_19_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_19_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_19_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_19_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_19_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_19_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_19_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_19_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_19_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_19_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_19_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_19_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_19_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_19_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_19_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_19_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_19_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_19_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_19_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_19_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_19_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_19_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_19_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_19_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_19_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_19_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_19_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_19_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_19_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_19_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_19_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_19_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_19_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_19_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_19_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_19_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_19_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_19_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_19_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_19_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_19_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_19_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_19_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_19_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_19_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_19_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_19_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_19_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_19_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_19_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_19_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_19_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_19_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_19_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_19_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N248, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N252, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N254, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N256, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N258, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N260, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N262, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N264, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N266, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N268, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N270, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N272, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N274, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N276, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N278, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N280, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N282, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N284, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N286, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N288, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N290, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N292, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N294, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N296, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N298, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N300, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N302, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N304, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N306, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N308, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N310, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N249, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N251, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N253, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N255, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N257, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N259, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N261, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N263, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N265, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N267, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N269, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N271, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N273, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N275, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N277, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N279, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N281, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N283, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N285, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N287, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N289, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N291, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N293, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N295, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N297, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N299, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N301, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N303, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N305, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N307, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N309, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N311, 
         -- Connections to port 'Z'
         Z(0) => N519 );
   C13072_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_18_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_18_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_18_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_18_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_18_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_18_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_18_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_18_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_18_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_18_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_18_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_18_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_18_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_18_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_18_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_18_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_18_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_18_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_18_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_18_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_18_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_18_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_18_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_18_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_18_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_18_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_18_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_18_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_18_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_18_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_18_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_18_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_18_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_18_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_18_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_18_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_18_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_18_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_18_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_18_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_18_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_18_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_18_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_18_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_18_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_18_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_18_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_18_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_18_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_18_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_18_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_18_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_18_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_18_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_18_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_18_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_18_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_18_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_18_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_18_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_18_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_18_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_18_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_18_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N248, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N252, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N254, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N256, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N258, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N260, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N262, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N264, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N266, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N268, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N270, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N272, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N274, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N276, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N278, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N280, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N282, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N284, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N286, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N288, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N290, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N292, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N294, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N296, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N298, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N300, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N302, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N304, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N306, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N308, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N310, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N249, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N251, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N253, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N255, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N257, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N259, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N261, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N263, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N265, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N267, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N269, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N271, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N273, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N275, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N277, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N279, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N281, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N283, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N285, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N287, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N289, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N291, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N293, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N295, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N297, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N299, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N301, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N303, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N305, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N307, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N309, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N311, 
         -- Connections to port 'Z'
         Z(0) => N520 );
   C13073_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_17_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_17_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_17_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_17_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_17_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_17_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_17_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_17_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_17_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_17_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_17_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_17_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_17_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_17_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_17_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_17_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_17_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_17_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_17_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_17_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_17_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_17_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_17_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_17_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_17_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_17_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_17_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_17_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_17_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_17_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_17_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_17_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_17_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_17_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_17_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_17_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_17_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_17_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_17_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_17_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_17_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_17_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_17_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_17_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_17_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_17_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_17_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_17_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_17_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_17_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_17_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_17_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_17_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_17_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_17_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_17_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_17_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_17_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_17_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_17_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_17_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_17_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_17_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_17_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N248, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N252, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N254, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N256, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N258, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N260, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N262, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N264, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N266, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N268, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N270, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N272, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N274, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N276, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N278, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N280, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N282, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N284, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N286, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N288, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N290, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N292, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N294, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N296, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N298, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N300, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N302, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N304, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N306, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N308, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N310, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N249, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N251, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N253, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N255, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N257, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N259, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N261, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N263, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N265, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N267, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N269, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N271, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N273, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N275, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N277, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N279, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N281, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N283, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N285, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N287, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N289, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N291, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N293, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N295, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N297, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N299, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N301, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N303, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N305, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N307, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N309, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N311, 
         -- Connections to port 'Z'
         Z(0) => N521 );
   C13074_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_16_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_16_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_16_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_16_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_16_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_16_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_16_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_16_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_16_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_16_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_16_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_16_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_16_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_16_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_16_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_16_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_16_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_16_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_16_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_16_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_16_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_16_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_16_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_16_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_16_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_16_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_16_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_16_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_16_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_16_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_16_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_16_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_16_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_16_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_16_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_16_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_16_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_16_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_16_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_16_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_16_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_16_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_16_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_16_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_16_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_16_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_16_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_16_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_16_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_16_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_16_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_16_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_16_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_16_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_16_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_16_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_16_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_16_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_16_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_16_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_16_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_16_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_16_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_16_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N248, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N252, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N254, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N256, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N258, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N260, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N262, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N264, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N266, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N268, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N270, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N272, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N274, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N276, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N278, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N280, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N282, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N284, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N286, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N288, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N290, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N292, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N294, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N296, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N298, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N300, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N302, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N304, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N306, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N308, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N310, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N249, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N251, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N253, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N255, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N257, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N259, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N261, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N263, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N265, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N267, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N269, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N271, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N273, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N275, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N277, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N279, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N281, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N283, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N285, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N287, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N289, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N291, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N293, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N295, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N297, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N299, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N301, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N303, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N305, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N307, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N309, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N311, 
         -- Connections to port 'Z'
         Z(0) => N522 );
   C13075_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_15_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_15_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_15_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_15_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_15_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_15_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_15_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_15_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_15_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_15_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_15_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_15_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_15_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_15_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_15_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_15_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_15_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_15_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_15_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_15_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_15_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_15_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_15_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_15_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_15_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_15_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_15_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_15_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_15_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_15_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_15_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_15_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_15_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_15_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_15_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_15_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_15_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_15_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_15_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_15_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_15_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_15_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_15_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_15_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_15_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_15_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_15_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_15_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_15_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_15_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_15_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_15_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_15_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_15_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_15_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_15_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_15_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_15_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_15_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_15_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_15_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_15_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_15_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_15_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N248, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N252, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N254, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N256, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N258, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N260, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N262, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N264, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N266, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N268, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N270, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N272, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N274, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N276, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N278, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N280, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N282, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N284, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N286, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N288, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N290, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N292, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N294, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N296, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N298, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N300, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N302, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N304, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N306, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N308, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N310, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N249, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N251, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N253, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N255, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N257, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N259, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N261, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N263, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N265, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N267, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N269, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N271, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N273, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N275, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N277, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N279, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N281, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N283, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N285, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N287, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N289, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N291, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N293, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N295, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N297, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N299, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N301, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N303, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N305, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N307, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N309, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N311, 
         -- Connections to port 'Z'
         Z(0) => N523 );
   C13076_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_14_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_14_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_14_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_14_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_14_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_14_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_14_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_14_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_14_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_14_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_14_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_14_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_14_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_14_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_14_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_14_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_14_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_14_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_14_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_14_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_14_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_14_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_14_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_14_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_14_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_14_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_14_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_14_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_14_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_14_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_14_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_14_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_14_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_14_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_14_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_14_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_14_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_14_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_14_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_14_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_14_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_14_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_14_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_14_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_14_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_14_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_14_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_14_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_14_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_14_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_14_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_14_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_14_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_14_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_14_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_14_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_14_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_14_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_14_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_14_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_14_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_14_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_14_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_14_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N248, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N252, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N254, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N256, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N258, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N260, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N262, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N264, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N266, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N268, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N270, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N272, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N274, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N276, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N278, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N280, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N282, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N284, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N286, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N288, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N290, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N292, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N294, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N296, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N298, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N300, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N302, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N304, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N306, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N308, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N310, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N249, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N251, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N253, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N255, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N257, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N259, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N261, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N263, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N265, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N267, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N269, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N271, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N273, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N275, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N277, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N279, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N281, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N283, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N285, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N287, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N289, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N291, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N293, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N295, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N297, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N299, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N301, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N303, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N305, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N307, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N309, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N311, 
         -- Connections to port 'Z'
         Z(0) => N524 );
   C13077_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_13_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_13_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_13_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_13_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_13_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_13_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_13_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_13_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_13_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_13_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_13_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_13_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_13_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_13_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_13_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_13_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_13_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_13_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_13_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_13_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_13_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_13_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_13_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_13_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_13_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_13_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_13_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_13_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_13_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_13_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_13_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_13_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_13_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_13_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_13_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_13_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_13_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_13_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_13_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_13_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_13_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_13_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_13_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_13_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_13_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_13_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_13_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_13_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_13_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_13_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_13_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_13_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_13_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_13_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_13_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_13_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_13_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_13_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_13_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_13_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_13_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_13_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_13_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_13_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N248, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N252, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N254, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N256, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N258, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N260, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N262, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N264, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N266, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N268, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N270, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N272, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N274, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N276, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N278, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N280, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N282, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N284, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N286, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N288, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N290, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N292, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N294, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N296, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N298, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N300, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N302, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N304, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N306, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N308, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N310, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N249, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N251, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N253, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N255, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N257, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N259, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N261, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N263, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N265, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N267, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N269, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N271, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N273, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N275, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N277, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N279, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N281, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N283, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N285, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N287, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N289, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N291, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N293, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N295, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N297, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N299, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N301, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N303, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N305, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N307, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N309, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N311, 
         -- Connections to port 'Z'
         Z(0) => N525 );
   C13078_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_12_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_12_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_12_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_12_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_12_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_12_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_12_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_12_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_12_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_12_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_12_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_12_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_12_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_12_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_12_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_12_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_12_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_12_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_12_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_12_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_12_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_12_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_12_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_12_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_12_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_12_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_12_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_12_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_12_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_12_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_12_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_12_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_12_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_12_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_12_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_12_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_12_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_12_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_12_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_12_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_12_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_12_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_12_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_12_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_12_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_12_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_12_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_12_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_12_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_12_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_12_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_12_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_12_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_12_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_12_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_12_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_12_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_12_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_12_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_12_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_12_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_12_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_12_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_12_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N248, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N252, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N254, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N256, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N258, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N260, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N262, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N264, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N266, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N268, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N270, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N272, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N274, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N276, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N278, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N280, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N282, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N284, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N286, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N288, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N290, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N292, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N294, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N296, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N298, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N300, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N302, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N304, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N306, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N308, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N310, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N249, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N251, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N253, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N255, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N257, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N259, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N261, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N263, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N265, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N267, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N269, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N271, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N273, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N275, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N277, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N279, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N281, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N283, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N285, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N287, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N289, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N291, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N293, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N295, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N297, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N299, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N301, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N303, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N305, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N307, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N309, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N311, 
         -- Connections to port 'Z'
         Z(0) => N526 );
   C13079_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_11_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_11_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_11_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_11_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_11_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_11_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_11_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_11_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_11_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_11_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_11_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_11_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_11_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_11_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_11_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_11_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_11_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_11_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_11_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_11_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_11_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_11_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_11_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_11_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_11_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_11_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_11_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_11_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_11_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_11_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_11_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_11_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_11_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_11_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_11_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_11_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_11_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_11_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_11_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_11_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_11_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_11_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_11_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_11_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_11_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_11_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_11_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_11_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_11_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_11_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_11_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_11_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_11_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_11_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_11_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_11_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_11_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_11_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_11_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_11_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_11_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_11_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_11_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_11_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N248, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N252, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N254, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N256, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N258, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N260, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N262, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N264, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N266, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N268, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N270, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N272, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N274, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N276, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N278, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N280, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N282, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N284, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N286, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N288, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N290, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N292, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N294, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N296, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N298, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N300, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N302, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N304, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N306, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N308, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N310, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N249, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N251, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N253, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N255, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N257, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N259, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N261, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N263, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N265, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N267, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N269, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N271, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N273, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N275, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N277, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N279, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N281, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N283, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N285, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N287, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N289, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N291, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N293, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N295, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N297, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N299, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N301, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N303, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N305, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N307, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N309, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N311, 
         -- Connections to port 'Z'
         Z(0) => N527 );
   C13080_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_10_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_10_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_10_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_10_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_10_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_10_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_10_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_10_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_10_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_10_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_10_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_10_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_10_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_10_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_10_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_10_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_10_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_10_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_10_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_10_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_10_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_10_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_10_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_10_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_10_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_10_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_10_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_10_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_10_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_10_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_10_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_10_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_10_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_10_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_10_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_10_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_10_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_10_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_10_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_10_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_10_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_10_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_10_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_10_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_10_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_10_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_10_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_10_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_10_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_10_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_10_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_10_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_10_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_10_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_10_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_10_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_10_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_10_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_10_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_10_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_10_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_10_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_10_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_10_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N248, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N252, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N254, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N256, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N258, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N260, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N262, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N264, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N266, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N268, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N270, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N272, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N274, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N276, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N278, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N280, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N282, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N284, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N286, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N288, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N290, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N292, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N294, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N296, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N298, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N300, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N302, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N304, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N306, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N308, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N310, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N249, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N251, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N253, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N255, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N257, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N259, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N261, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N263, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N265, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N267, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N269, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N271, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N273, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N275, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N277, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N279, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N281, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N283, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N285, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N287, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N289, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N291, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N293, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N295, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N297, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N299, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N301, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N303, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N305, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N307, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N309, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N311, 
         -- Connections to port 'Z'
         Z(0) => N528 );
   C13081_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_9_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_9_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_9_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_9_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_9_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_9_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_9_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_9_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_9_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_9_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_9_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_9_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_9_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_9_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_9_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_9_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_9_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_9_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_9_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_9_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_9_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_9_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_9_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_9_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_9_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_9_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_9_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_9_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_9_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_9_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_9_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_9_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_9_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_9_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_9_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_9_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_9_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_9_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_9_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_9_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_9_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_9_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_9_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_9_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_9_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_9_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_9_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_9_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_9_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_9_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_9_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_9_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_9_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_9_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_9_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_9_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_9_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_9_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_9_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_9_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_9_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_9_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_9_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_9_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N248, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N252, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N254, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N256, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N258, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N260, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N262, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N264, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N266, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N268, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N270, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N272, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N274, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N276, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N278, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N280, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N282, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N284, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N286, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N288, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N290, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N292, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N294, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N296, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N298, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N300, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N302, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N304, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N306, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N308, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N310, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N249, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N251, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N253, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N255, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N257, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N259, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N261, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N263, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N265, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N267, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N269, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N271, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N273, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N275, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N277, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N279, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N281, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N283, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N285, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N287, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N289, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N291, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N293, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N295, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N297, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N299, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N301, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N303, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N305, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N307, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N309, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N311, 
         -- Connections to port 'Z'
         Z(0) => N529 );
   C13082_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_8_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_8_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_8_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_8_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_8_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_8_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_8_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_8_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_8_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_8_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_8_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_8_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_8_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_8_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_8_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_8_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_8_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_8_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_8_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_8_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_8_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_8_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_8_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_8_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_8_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_8_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_8_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_8_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_8_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_8_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_8_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_8_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_8_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_8_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_8_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_8_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_8_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_8_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_8_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_8_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_8_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_8_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_8_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_8_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_8_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_8_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_8_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_8_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_8_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_8_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_8_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_8_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_8_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_8_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_8_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_8_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_8_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_8_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_8_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_8_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_8_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_8_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_8_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_8_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N248, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N252, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N254, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N256, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N258, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N260, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N262, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N264, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N266, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N268, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N270, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N272, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N274, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N276, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N278, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N280, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N282, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N284, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N286, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N288, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N290, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N292, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N294, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N296, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N298, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N300, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N302, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N304, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N306, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N308, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N310, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N249, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N251, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N253, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N255, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N257, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N259, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N261, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N263, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N265, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N267, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N269, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N271, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N273, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N275, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N277, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N279, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N281, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N283, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N285, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N287, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N289, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N291, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N293, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N295, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N297, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N299, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N301, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N303, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N305, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N307, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N309, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N311, 
         -- Connections to port 'Z'
         Z(0) => N530 );
   C13083_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_7_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_7_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_7_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_7_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_7_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_7_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_7_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_7_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_7_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_7_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_7_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_7_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_7_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_7_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_7_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_7_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_7_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_7_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_7_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_7_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_7_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_7_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_7_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_7_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_7_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_7_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_7_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_7_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_7_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_7_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_7_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_7_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_7_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_7_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_7_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_7_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_7_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_7_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_7_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_7_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_7_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_7_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_7_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_7_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_7_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_7_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_7_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_7_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_7_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_7_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_7_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_7_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_7_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_7_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_7_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_7_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_7_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_7_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_7_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_7_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_7_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_7_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_7_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_7_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N248, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N252, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N254, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N256, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N258, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N260, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N262, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N264, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N266, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N268, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N270, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N272, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N274, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N276, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N278, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N280, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N282, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N284, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N286, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N288, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N290, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N292, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N294, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N296, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N298, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N300, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N302, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N304, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N306, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N308, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N310, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N249, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N251, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N253, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N255, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N257, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N259, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N261, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N263, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N265, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N267, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N269, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N271, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N273, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N275, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N277, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N279, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N281, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N283, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N285, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N287, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N289, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N291, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N293, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N295, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N297, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N299, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N301, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N303, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N305, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N307, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N309, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N311, 
         -- Connections to port 'Z'
         Z(0) => N531 );
   C13084_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_6_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_6_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_6_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_6_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_6_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_6_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_6_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_6_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_6_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_6_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_6_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_6_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_6_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_6_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_6_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_6_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_6_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_6_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_6_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_6_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_6_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_6_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_6_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_6_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_6_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_6_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_6_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_6_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_6_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_6_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_6_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_6_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_6_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_6_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_6_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_6_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_6_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_6_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_6_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_6_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_6_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_6_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_6_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_6_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_6_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_6_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_6_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_6_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_6_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_6_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_6_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_6_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_6_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_6_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_6_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_6_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_6_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_6_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_6_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_6_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_6_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_6_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_6_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_6_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N248, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N252, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N254, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N256, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N258, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N260, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N262, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N264, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N266, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N268, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N270, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N272, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N274, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N276, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N278, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N280, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N282, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N284, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N286, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N288, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N290, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N292, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N294, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N296, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N298, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N300, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N302, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N304, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N306, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N308, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N310, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N249, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N251, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N253, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N255, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N257, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N259, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N261, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N263, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N265, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N267, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N269, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N271, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N273, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N275, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N277, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N279, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N281, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N283, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N285, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N287, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N289, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N291, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N293, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N295, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N297, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N299, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N301, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N303, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N305, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N307, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N309, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N311, 
         -- Connections to port 'Z'
         Z(0) => N532 );
   C13085_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_5_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_5_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_5_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_5_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_5_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_5_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_5_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_5_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_5_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_5_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_5_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_5_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_5_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_5_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_5_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_5_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_5_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_5_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_5_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_5_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_5_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_5_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_5_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_5_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_5_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_5_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_5_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_5_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_5_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_5_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_5_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_5_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_5_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_5_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_5_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_5_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_5_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_5_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_5_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_5_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_5_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_5_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_5_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_5_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_5_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_5_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_5_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_5_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_5_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_5_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_5_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_5_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_5_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_5_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_5_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_5_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_5_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_5_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_5_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_5_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_5_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_5_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_5_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_5_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N248, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N252, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N254, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N256, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N258, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N260, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N262, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N264, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N266, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N268, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N270, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N272, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N274, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N276, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N278, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N280, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N282, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N284, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N286, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N288, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N290, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N292, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N294, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N296, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N298, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N300, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N302, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N304, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N306, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N308, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N310, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N249, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N251, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N253, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N255, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N257, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N259, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N261, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N263, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N265, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N267, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N269, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N271, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N273, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N275, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N277, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N279, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N281, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N283, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N285, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N287, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N289, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N291, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N293, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N295, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N297, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N299, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N301, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N303, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N305, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N307, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N309, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N311, 
         -- Connections to port 'Z'
         Z(0) => N533 );
   C13086_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_4_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_4_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_4_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_4_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_4_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_4_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_4_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_4_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_4_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_4_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_4_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_4_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_4_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_4_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_4_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_4_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_4_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_4_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_4_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_4_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_4_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_4_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_4_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_4_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_4_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_4_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_4_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_4_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_4_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_4_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_4_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_4_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_4_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_4_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_4_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_4_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_4_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_4_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_4_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_4_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_4_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_4_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_4_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_4_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_4_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_4_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_4_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_4_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_4_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_4_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_4_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_4_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_4_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_4_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_4_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_4_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_4_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_4_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_4_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_4_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_4_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_4_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_4_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_4_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N248, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N252, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N254, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N256, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N258, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N260, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N262, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N264, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N266, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N268, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N270, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N272, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N274, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N276, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N278, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N280, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N282, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N284, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N286, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N288, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N290, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N292, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N294, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N296, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N298, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N300, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N302, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N304, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N306, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N308, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N310, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N249, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N251, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N253, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N255, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N257, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N259, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N261, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N263, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N265, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N267, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N269, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N271, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N273, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N275, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N277, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N279, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N281, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N283, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N285, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N287, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N289, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N291, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N293, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N295, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N297, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N299, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N301, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N303, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N305, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N307, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N309, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N311, 
         -- Connections to port 'Z'
         Z(0) => N534 );
   C13087_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_3_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_3_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_3_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_3_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_3_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_3_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_3_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_3_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_3_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_3_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_3_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_3_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_3_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_3_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_3_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_3_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_3_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_3_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_3_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_3_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_3_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_3_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_3_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_3_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_3_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_3_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_3_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_3_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_3_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_3_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_3_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_3_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_3_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_3_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_3_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_3_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_3_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_3_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_3_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_3_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_3_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_3_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_3_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_3_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_3_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_3_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_3_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_3_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_3_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_3_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_3_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_3_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_3_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_3_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_3_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_3_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_3_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_3_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_3_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_3_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_3_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_3_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_3_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_3_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N248, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N252, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N254, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N256, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N258, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N260, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N262, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N264, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N266, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N268, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N270, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N272, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N274, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N276, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N278, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N280, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N282, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N284, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N286, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N288, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N290, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N292, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N294, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N296, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N298, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N300, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N302, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N304, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N306, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N308, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N310, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N249, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N251, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N253, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N255, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N257, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N259, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N261, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N263, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N265, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N267, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N269, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N271, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N273, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N275, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N277, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N279, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N281, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N283, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N285, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N287, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N289, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N291, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N293, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N295, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N297, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N299, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N301, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N303, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N305, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N307, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N309, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N311, 
         -- Connections to port 'Z'
         Z(0) => N535 );
   C13088_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_2_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_2_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_2_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_2_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_2_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_2_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_2_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_2_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_2_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_2_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_2_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_2_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_2_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_2_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_2_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_2_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_2_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_2_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_2_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_2_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_2_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_2_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_2_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_2_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_2_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_2_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_2_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_2_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_2_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_2_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_2_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_2_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_2_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_2_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_2_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_2_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_2_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_2_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_2_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_2_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_2_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_2_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_2_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_2_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_2_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_2_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_2_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_2_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_2_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_2_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_2_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_2_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_2_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_2_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_2_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_2_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_2_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_2_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_2_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_2_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_2_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_2_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_2_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_2_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N248, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N252, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N254, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N256, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N258, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N260, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N262, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N264, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N266, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N268, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N270, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N272, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N274, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N276, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N278, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N280, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N282, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N284, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N286, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N288, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N290, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N292, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N294, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N296, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N298, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N300, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N302, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N304, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N306, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N308, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N310, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N249, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N251, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N253, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N255, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N257, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N259, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N261, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N263, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N265, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N267, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N269, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N271, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N273, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N275, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N277, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N279, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N281, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N283, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N285, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N287, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N289, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N291, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N293, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N295, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N297, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N299, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N301, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N303, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N305, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N307, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N309, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N311, 
         -- Connections to port 'Z'
         Z(0) => N536 );
   C13089_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_1_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_1_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_1_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_1_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_1_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_1_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_1_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_1_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_1_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_1_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_1_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_1_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_1_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_1_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_1_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_1_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_1_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_1_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_1_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_1_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_1_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_1_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_1_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_1_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_1_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_1_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_1_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_1_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_1_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_1_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_1_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_1_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_1_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_1_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_1_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_1_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_1_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_1_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_1_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_1_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_1_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_1_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_1_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_1_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_1_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_1_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_1_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_1_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_1_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_1_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_1_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_1_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_1_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_1_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_1_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_1_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_1_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_1_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_1_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_1_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_1_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_1_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_1_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_1_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N248, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N252, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N254, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N256, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N258, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N260, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N262, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N264, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N266, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N268, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N270, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N272, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N274, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N276, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N278, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N280, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N282, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N284, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N286, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N288, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N290, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N292, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N294, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N296, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N298, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N300, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N302, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N304, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N306, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N308, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N310, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N249, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N251, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N253, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N255, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N257, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N259, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N261, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N263, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N265, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N267, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N269, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N271, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N273, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N275, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N277, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N279, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N281, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N283, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N285, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N287, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N289, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N291, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N293, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N295, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N297, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N299, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N301, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N303, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N305, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N307, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N309, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N311, 
         -- Connections to port 'Z'
         Z(0) => N537 );
   C13090_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_0_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_0_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_0_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_0_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_0_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_0_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_0_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_0_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_0_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_0_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_0_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_0_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_0_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_0_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_0_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_0_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_0_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_0_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_0_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_0_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_0_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_0_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_0_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_0_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_0_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_0_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_0_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_0_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_0_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_0_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_0_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_0_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_0_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_0_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_0_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_0_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_0_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_0_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_0_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_0_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_0_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_0_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_0_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_0_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_0_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_0_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_0_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_0_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_0_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_0_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_0_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_0_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_0_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_0_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_0_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_0_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_0_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_0_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_0_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_0_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_0_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_0_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N248, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N252, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N254, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N256, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N258, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N260, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N262, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N264, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N266, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N268, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N270, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N272, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N274, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N276, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N278, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N280, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N282, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N284, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N286, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N288, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N290, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N292, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N294, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N296, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N298, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N300, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N302, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N304, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N306, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N308, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N310, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N249, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N251, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N253, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N255, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N257, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N259, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N261, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N263, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N265, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N267, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N269, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N271, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N273, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N275, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N277, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N279, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N281, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N283, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N285, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N287, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N289, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N291, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N293, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N295, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N297, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N299, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N301, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N303, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N305, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N307, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N309, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N311, 
         -- Connections to port 'Z'
         Z(0) => N538 );
   C13227_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_31_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_31_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_31_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_31_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_31_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_31_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_31_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_31_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_31_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_31_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_31_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_31_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_31_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_31_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_31_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_31_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_31_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_31_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_31_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_31_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_31_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_31_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_31_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_31_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_31_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_31_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_31_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_31_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_31_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_31_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_31_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_31_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_31_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_31_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_31_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_31_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_31_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_31_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_31_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_31_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_31_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_31_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_31_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_31_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_31_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_31_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_31_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_31_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_31_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_31_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_31_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_31_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_31_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_31_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_31_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_31_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_31_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_31_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_31_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_31_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_31_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_31_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_31_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_31_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N410, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N412, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N414, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N416, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N418, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N420, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N422, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N424, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N426, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N428, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N430, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N432, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N434, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N436, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N438, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N440, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N442, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N444, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N446, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N448, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N450, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N452, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N454, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N456, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N458, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N460, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N462, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N464, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N466, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N468, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N470, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N472, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N411, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N413, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N415, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N417, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N419, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N421, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N423, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N425, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N427, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N429, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N431, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N433, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N435, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N437, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N439, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N441, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N443, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N445, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N447, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N449, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N451, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N453, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N455, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N457, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N459, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N461, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N463, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N465, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N467, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N469, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N471, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N473, 
         -- Connections to port 'Z'
         Z(0) => N539 );
   C13228_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_30_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_30_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_30_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_30_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_30_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_30_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_30_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_30_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_30_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_30_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_30_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_30_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_30_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_30_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_30_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_30_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_30_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_30_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_30_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_30_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_30_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_30_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_30_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_30_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_30_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_30_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_30_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_30_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_30_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_30_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_30_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_30_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_30_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_30_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_30_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_30_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_30_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_30_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_30_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_30_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_30_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_30_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_30_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_30_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_30_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_30_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_30_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_30_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_30_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_30_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_30_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_30_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_30_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_30_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_30_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_30_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_30_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_30_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_30_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_30_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_30_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_30_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_30_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_30_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N410, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N412, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N414, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N416, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N418, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N420, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N422, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N424, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N426, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N428, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N430, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N432, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N434, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N436, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N438, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N440, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N442, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N444, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N446, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N448, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N450, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N452, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N454, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N456, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N458, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N460, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N462, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N464, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N466, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N468, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N470, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N472, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N411, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N413, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N415, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N417, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N419, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N421, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N423, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N425, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N427, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N429, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N431, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N433, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N435, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N437, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N439, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N441, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N443, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N445, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N447, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N449, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N451, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N453, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N455, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N457, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N459, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N461, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N463, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N465, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N467, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N469, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N471, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N473, 
         -- Connections to port 'Z'
         Z(0) => N540 );
   C13229_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_29_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_29_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_29_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_29_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_29_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_29_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_29_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_29_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_29_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_29_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_29_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_29_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_29_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_29_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_29_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_29_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_29_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_29_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_29_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_29_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_29_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_29_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_29_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_29_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_29_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_29_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_29_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_29_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_29_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_29_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_29_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_29_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_29_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_29_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_29_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_29_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_29_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_29_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_29_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_29_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_29_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_29_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_29_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_29_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_29_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_29_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_29_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_29_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_29_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_29_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_29_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_29_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_29_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_29_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_29_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_29_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_29_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_29_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_29_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_29_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_29_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_29_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_29_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_29_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N410, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N412, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N414, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N416, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N418, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N420, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N422, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N424, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N426, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N428, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N430, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N432, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N434, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N436, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N438, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N440, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N442, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N444, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N446, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N448, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N450, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N452, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N454, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N456, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N458, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N460, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N462, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N464, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N466, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N468, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N470, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N472, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N411, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N413, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N415, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N417, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N419, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N421, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N423, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N425, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N427, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N429, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N431, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N433, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N435, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N437, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N439, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N441, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N443, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N445, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N447, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N449, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N451, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N453, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N455, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N457, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N459, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N461, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N463, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N465, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N467, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N469, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N471, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N473, 
         -- Connections to port 'Z'
         Z(0) => N541 );
   C13230_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_28_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_28_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_28_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_28_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_28_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_28_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_28_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_28_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_28_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_28_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_28_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_28_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_28_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_28_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_28_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_28_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_28_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_28_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_28_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_28_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_28_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_28_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_28_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_28_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_28_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_28_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_28_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_28_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_28_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_28_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_28_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_28_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_28_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_28_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_28_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_28_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_28_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_28_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_28_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_28_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_28_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_28_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_28_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_28_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_28_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_28_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_28_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_28_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_28_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_28_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_28_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_28_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_28_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_28_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_28_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_28_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_28_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_28_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_28_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_28_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_28_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_28_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_28_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_28_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N410, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N412, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N414, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N416, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N418, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N420, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N422, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N424, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N426, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N428, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N430, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N432, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N434, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N436, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N438, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N440, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N442, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N444, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N446, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N448, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N450, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N452, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N454, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N456, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N458, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N460, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N462, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N464, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N466, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N468, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N470, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N472, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N411, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N413, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N415, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N417, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N419, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N421, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N423, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N425, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N427, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N429, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N431, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N433, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N435, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N437, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N439, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N441, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N443, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N445, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N447, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N449, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N451, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N453, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N455, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N457, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N459, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N461, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N463, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N465, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N467, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N469, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N471, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N473, 
         -- Connections to port 'Z'
         Z(0) => N542 );
   C13231_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_27_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_27_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_27_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_27_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_27_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_27_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_27_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_27_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_27_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_27_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_27_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_27_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_27_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_27_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_27_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_27_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_27_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_27_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_27_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_27_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_27_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_27_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_27_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_27_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_27_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_27_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_27_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_27_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_27_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_27_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_27_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_27_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_27_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_27_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_27_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_27_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_27_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_27_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_27_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_27_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_27_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_27_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_27_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_27_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_27_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_27_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_27_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_27_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_27_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_27_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_27_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_27_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_27_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_27_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_27_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_27_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_27_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_27_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_27_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_27_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_27_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_27_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_27_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_27_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N410, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N412, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N414, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N416, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N418, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N420, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N422, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N424, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N426, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N428, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N430, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N432, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N434, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N436, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N438, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N440, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N442, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N444, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N446, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N448, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N450, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N452, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N454, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N456, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N458, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N460, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N462, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N464, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N466, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N468, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N470, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N472, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N411, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N413, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N415, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N417, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N419, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N421, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N423, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N425, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N427, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N429, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N431, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N433, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N435, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N437, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N439, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N441, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N443, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N445, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N447, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N449, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N451, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N453, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N455, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N457, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N459, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N461, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N463, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N465, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N467, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N469, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N471, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N473, 
         -- Connections to port 'Z'
         Z(0) => N543 );
   C13232_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_26_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_26_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_26_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_26_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_26_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_26_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_26_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_26_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_26_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_26_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_26_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_26_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_26_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_26_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_26_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_26_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_26_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_26_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_26_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_26_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_26_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_26_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_26_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_26_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_26_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_26_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_26_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_26_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_26_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_26_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_26_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_26_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_26_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_26_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_26_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_26_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_26_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_26_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_26_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_26_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_26_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_26_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_26_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_26_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_26_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_26_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_26_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_26_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_26_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_26_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_26_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_26_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_26_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_26_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_26_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_26_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_26_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_26_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_26_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_26_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_26_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_26_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_26_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_26_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N410, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N412, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N414, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N416, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N418, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N420, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N422, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N424, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N426, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N428, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N430, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N432, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N434, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N436, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N438, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N440, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N442, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N444, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N446, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N448, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N450, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N452, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N454, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N456, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N458, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N460, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N462, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N464, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N466, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N468, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N470, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N472, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N411, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N413, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N415, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N417, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N419, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N421, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N423, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N425, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N427, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N429, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N431, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N433, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N435, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N437, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N439, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N441, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N443, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N445, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N447, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N449, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N451, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N453, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N455, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N457, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N459, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N461, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N463, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N465, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N467, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N469, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N471, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N473, 
         -- Connections to port 'Z'
         Z(0) => N544 );
   C13233_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_25_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_25_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_25_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_25_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_25_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_25_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_25_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_25_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_25_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_25_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_25_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_25_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_25_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_25_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_25_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_25_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_25_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_25_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_25_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_25_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_25_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_25_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_25_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_25_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_25_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_25_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_25_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_25_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_25_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_25_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_25_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_25_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_25_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_25_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_25_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_25_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_25_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_25_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_25_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_25_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_25_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_25_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_25_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_25_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_25_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_25_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_25_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_25_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_25_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_25_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_25_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_25_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_25_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_25_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_25_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_25_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_25_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_25_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_25_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_25_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_25_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_25_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_25_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_25_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N410, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N412, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N414, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N416, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N418, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N420, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N422, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N424, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N426, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N428, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N430, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N432, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N434, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N436, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N438, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N440, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N442, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N444, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N446, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N448, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N450, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N452, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N454, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N456, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N458, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N460, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N462, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N464, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N466, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N468, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N470, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N472, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N411, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N413, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N415, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N417, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N419, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N421, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N423, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N425, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N427, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N429, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N431, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N433, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N435, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N437, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N439, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N441, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N443, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N445, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N447, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N449, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N451, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N453, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N455, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N457, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N459, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N461, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N463, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N465, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N467, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N469, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N471, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N473, 
         -- Connections to port 'Z'
         Z(0) => N545 );
   C13234_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_24_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_24_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_24_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_24_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_24_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_24_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_24_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_24_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_24_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_24_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_24_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_24_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_24_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_24_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_24_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_24_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_24_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_24_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_24_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_24_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_24_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_24_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_24_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_24_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_24_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_24_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_24_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_24_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_24_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_24_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_24_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_24_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_24_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_24_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_24_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_24_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_24_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_24_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_24_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_24_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_24_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_24_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_24_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_24_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_24_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_24_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_24_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_24_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_24_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_24_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_24_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_24_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_24_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_24_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_24_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_24_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_24_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_24_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_24_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_24_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_24_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_24_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_24_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_24_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N410, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N412, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N414, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N416, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N418, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N420, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N422, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N424, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N426, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N428, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N430, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N432, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N434, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N436, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N438, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N440, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N442, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N444, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N446, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N448, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N450, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N452, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N454, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N456, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N458, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N460, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N462, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N464, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N466, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N468, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N470, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N472, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N411, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N413, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N415, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N417, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N419, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N421, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N423, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N425, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N427, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N429, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N431, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N433, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N435, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N437, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N439, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N441, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N443, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N445, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N447, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N449, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N451, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N453, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N455, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N457, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N459, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N461, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N463, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N465, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N467, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N469, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N471, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N473, 
         -- Connections to port 'Z'
         Z(0) => N546 );
   C13235_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_23_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_23_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_23_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_23_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_23_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_23_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_23_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_23_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_23_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_23_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_23_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_23_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_23_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_23_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_23_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_23_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_23_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_23_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_23_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_23_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_23_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_23_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_23_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_23_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_23_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_23_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_23_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_23_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_23_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_23_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_23_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_23_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_23_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_23_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_23_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_23_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_23_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_23_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_23_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_23_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_23_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_23_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_23_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_23_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_23_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_23_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_23_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_23_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_23_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_23_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_23_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_23_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_23_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_23_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_23_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_23_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_23_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_23_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_23_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_23_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_23_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_23_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_23_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_23_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N410, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N412, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N414, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N416, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N418, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N420, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N422, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N424, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N426, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N428, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N430, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N432, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N434, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N436, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N438, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N440, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N442, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N444, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N446, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N448, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N450, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N452, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N454, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N456, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N458, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N460, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N462, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N464, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N466, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N468, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N470, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N472, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N411, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N413, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N415, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N417, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N419, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N421, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N423, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N425, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N427, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N429, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N431, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N433, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N435, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N437, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N439, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N441, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N443, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N445, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N447, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N449, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N451, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N453, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N455, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N457, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N459, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N461, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N463, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N465, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N467, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N469, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N471, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N473, 
         -- Connections to port 'Z'
         Z(0) => N547 );
   C13236_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_22_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_22_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_22_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_22_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_22_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_22_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_22_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_22_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_22_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_22_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_22_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_22_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_22_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_22_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_22_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_22_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_22_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_22_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_22_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_22_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_22_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_22_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_22_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_22_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_22_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_22_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_22_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_22_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_22_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_22_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_22_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_22_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_22_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_22_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_22_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_22_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_22_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_22_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_22_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_22_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_22_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_22_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_22_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_22_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_22_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_22_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_22_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_22_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_22_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_22_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_22_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_22_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_22_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_22_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_22_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_22_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_22_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_22_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_22_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_22_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_22_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_22_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_22_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_22_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N410, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N412, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N414, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N416, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N418, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N420, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N422, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N424, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N426, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N428, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N430, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N432, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N434, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N436, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N438, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N440, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N442, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N444, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N446, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N448, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N450, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N452, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N454, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N456, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N458, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N460, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N462, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N464, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N466, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N468, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N470, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N472, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N411, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N413, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N415, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N417, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N419, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N421, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N423, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N425, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N427, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N429, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N431, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N433, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N435, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N437, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N439, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N441, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N443, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N445, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N447, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N449, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N451, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N453, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N455, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N457, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N459, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N461, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N463, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N465, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N467, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N469, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N471, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N473, 
         -- Connections to port 'Z'
         Z(0) => N548 );
   C13237_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_21_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_21_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_21_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_21_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_21_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_21_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_21_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_21_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_21_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_21_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_21_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_21_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_21_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_21_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_21_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_21_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_21_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_21_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_21_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_21_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_21_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_21_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_21_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_21_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_21_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_21_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_21_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_21_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_21_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_21_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_21_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_21_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_21_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_21_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_21_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_21_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_21_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_21_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_21_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_21_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_21_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_21_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_21_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_21_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_21_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_21_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_21_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_21_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_21_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_21_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_21_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_21_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_21_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_21_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_21_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_21_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_21_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_21_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_21_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_21_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_21_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_21_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_21_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_21_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N410, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N412, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N414, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N416, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N418, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N420, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N422, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N424, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N426, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N428, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N430, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N432, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N434, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N436, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N438, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N440, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N442, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N444, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N446, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N448, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N450, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N452, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N454, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N456, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N458, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N460, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N462, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N464, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N466, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N468, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N470, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N472, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N411, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N413, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N415, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N417, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N419, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N421, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N423, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N425, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N427, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N429, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N431, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N433, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N435, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N437, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N439, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N441, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N443, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N445, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N447, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N449, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N451, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N453, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N455, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N457, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N459, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N461, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N463, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N465, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N467, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N469, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N471, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N473, 
         -- Connections to port 'Z'
         Z(0) => N549 );
   C13238_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_20_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_20_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_20_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_20_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_20_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_20_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_20_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_20_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_20_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_20_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_20_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_20_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_20_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_20_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_20_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_20_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_20_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_20_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_20_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_20_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_20_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_20_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_20_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_20_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_20_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_20_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_20_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_20_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_20_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_20_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_20_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_20_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_20_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_20_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_20_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_20_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_20_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_20_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_20_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_20_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_20_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_20_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_20_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_20_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_20_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_20_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_20_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_20_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_20_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_20_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_20_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_20_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_20_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_20_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_20_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_20_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_20_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_20_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_20_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_20_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_20_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_20_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_20_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_20_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N410, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N412, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N414, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N416, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N418, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N420, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N422, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N424, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N426, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N428, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N430, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N432, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N434, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N436, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N438, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N440, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N442, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N444, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N446, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N448, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N450, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N452, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N454, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N456, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N458, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N460, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N462, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N464, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N466, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N468, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N470, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N472, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N411, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N413, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N415, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N417, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N419, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N421, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N423, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N425, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N427, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N429, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N431, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N433, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N435, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N437, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N439, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N441, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N443, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N445, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N447, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N449, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N451, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N453, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N455, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N457, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N459, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N461, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N463, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N465, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N467, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N469, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N471, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N473, 
         -- Connections to port 'Z'
         Z(0) => N550 );
   C13239_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_19_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_19_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_19_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_19_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_19_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_19_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_19_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_19_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_19_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_19_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_19_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_19_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_19_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_19_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_19_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_19_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_19_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_19_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_19_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_19_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_19_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_19_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_19_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_19_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_19_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_19_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_19_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_19_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_19_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_19_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_19_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_19_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_19_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_19_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_19_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_19_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_19_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_19_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_19_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_19_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_19_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_19_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_19_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_19_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_19_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_19_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_19_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_19_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_19_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_19_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_19_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_19_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_19_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_19_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_19_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_19_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_19_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_19_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_19_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_19_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_19_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_19_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_19_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_19_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N410, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N412, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N414, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N416, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N418, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N420, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N422, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N424, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N426, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N428, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N430, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N432, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N434, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N436, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N438, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N440, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N442, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N444, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N446, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N448, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N450, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N452, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N454, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N456, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N458, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N460, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N462, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N464, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N466, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N468, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N470, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N472, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N411, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N413, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N415, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N417, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N419, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N421, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N423, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N425, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N427, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N429, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N431, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N433, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N435, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N437, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N439, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N441, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N443, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N445, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N447, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N449, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N451, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N453, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N455, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N457, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N459, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N461, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N463, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N465, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N467, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N469, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N471, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N473, 
         -- Connections to port 'Z'
         Z(0) => N551 );
   C13240_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_18_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_18_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_18_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_18_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_18_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_18_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_18_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_18_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_18_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_18_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_18_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_18_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_18_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_18_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_18_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_18_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_18_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_18_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_18_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_18_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_18_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_18_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_18_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_18_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_18_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_18_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_18_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_18_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_18_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_18_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_18_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_18_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_18_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_18_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_18_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_18_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_18_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_18_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_18_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_18_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_18_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_18_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_18_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_18_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_18_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_18_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_18_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_18_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_18_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_18_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_18_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_18_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_18_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_18_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_18_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_18_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_18_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_18_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_18_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_18_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_18_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_18_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_18_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_18_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N410, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N412, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N414, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N416, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N418, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N420, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N422, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N424, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N426, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N428, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N430, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N432, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N434, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N436, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N438, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N440, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N442, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N444, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N446, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N448, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N450, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N452, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N454, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N456, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N458, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N460, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N462, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N464, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N466, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N468, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N470, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N472, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N411, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N413, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N415, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N417, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N419, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N421, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N423, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N425, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N427, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N429, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N431, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N433, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N435, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N437, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N439, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N441, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N443, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N445, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N447, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N449, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N451, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N453, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N455, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N457, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N459, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N461, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N463, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N465, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N467, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N469, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N471, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N473, 
         -- Connections to port 'Z'
         Z(0) => N552 );
   C13241_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_17_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_17_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_17_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_17_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_17_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_17_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_17_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_17_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_17_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_17_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_17_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_17_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_17_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_17_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_17_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_17_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_17_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_17_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_17_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_17_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_17_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_17_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_17_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_17_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_17_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_17_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_17_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_17_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_17_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_17_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_17_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_17_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_17_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_17_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_17_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_17_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_17_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_17_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_17_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_17_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_17_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_17_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_17_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_17_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_17_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_17_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_17_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_17_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_17_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_17_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_17_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_17_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_17_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_17_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_17_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_17_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_17_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_17_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_17_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_17_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_17_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_17_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_17_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_17_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N410, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N412, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N414, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N416, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N418, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N420, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N422, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N424, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N426, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N428, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N430, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N432, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N434, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N436, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N438, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N440, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N442, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N444, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N446, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N448, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N450, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N452, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N454, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N456, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N458, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N460, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N462, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N464, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N466, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N468, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N470, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N472, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N411, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N413, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N415, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N417, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N419, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N421, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N423, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N425, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N427, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N429, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N431, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N433, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N435, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N437, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N439, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N441, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N443, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N445, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N447, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N449, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N451, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N453, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N455, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N457, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N459, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N461, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N463, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N465, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N467, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N469, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N471, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N473, 
         -- Connections to port 'Z'
         Z(0) => N553 );
   C13242_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_16_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_16_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_16_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_16_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_16_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_16_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_16_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_16_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_16_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_16_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_16_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_16_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_16_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_16_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_16_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_16_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_16_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_16_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_16_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_16_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_16_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_16_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_16_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_16_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_16_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_16_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_16_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_16_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_16_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_16_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_16_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_16_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_16_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_16_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_16_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_16_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_16_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_16_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_16_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_16_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_16_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_16_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_16_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_16_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_16_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_16_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_16_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_16_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_16_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_16_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_16_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_16_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_16_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_16_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_16_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_16_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_16_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_16_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_16_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_16_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_16_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_16_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_16_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_16_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N410, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N412, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N414, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N416, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N418, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N420, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N422, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N424, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N426, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N428, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N430, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N432, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N434, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N436, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N438, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N440, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N442, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N444, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N446, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N448, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N450, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N452, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N454, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N456, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N458, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N460, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N462, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N464, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N466, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N468, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N470, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N472, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N411, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N413, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N415, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N417, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N419, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N421, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N423, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N425, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N427, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N429, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N431, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N433, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N435, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N437, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N439, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N441, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N443, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N445, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N447, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N449, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N451, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N453, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N455, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N457, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N459, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N461, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N463, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N465, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N467, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N469, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N471, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N473, 
         -- Connections to port 'Z'
         Z(0) => N554 );
   C13243_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_15_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_15_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_15_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_15_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_15_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_15_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_15_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_15_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_15_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_15_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_15_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_15_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_15_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_15_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_15_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_15_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_15_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_15_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_15_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_15_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_15_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_15_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_15_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_15_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_15_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_15_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_15_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_15_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_15_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_15_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_15_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_15_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_15_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_15_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_15_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_15_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_15_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_15_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_15_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_15_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_15_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_15_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_15_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_15_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_15_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_15_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_15_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_15_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_15_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_15_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_15_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_15_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_15_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_15_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_15_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_15_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_15_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_15_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_15_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_15_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_15_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_15_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_15_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_15_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N410, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N412, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N414, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N416, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N418, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N420, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N422, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N424, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N426, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N428, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N430, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N432, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N434, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N436, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N438, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N440, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N442, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N444, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N446, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N448, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N450, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N452, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N454, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N456, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N458, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N460, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N462, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N464, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N466, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N468, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N470, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N472, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N411, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N413, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N415, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N417, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N419, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N421, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N423, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N425, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N427, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N429, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N431, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N433, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N435, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N437, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N439, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N441, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N443, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N445, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N447, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N449, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N451, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N453, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N455, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N457, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N459, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N461, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N463, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N465, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N467, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N469, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N471, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N473, 
         -- Connections to port 'Z'
         Z(0) => N555 );
   C13244_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_14_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_14_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_14_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_14_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_14_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_14_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_14_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_14_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_14_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_14_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_14_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_14_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_14_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_14_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_14_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_14_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_14_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_14_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_14_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_14_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_14_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_14_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_14_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_14_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_14_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_14_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_14_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_14_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_14_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_14_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_14_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_14_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_14_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_14_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_14_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_14_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_14_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_14_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_14_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_14_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_14_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_14_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_14_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_14_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_14_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_14_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_14_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_14_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_14_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_14_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_14_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_14_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_14_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_14_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_14_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_14_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_14_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_14_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_14_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_14_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_14_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_14_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_14_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_14_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N410, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N412, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N414, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N416, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N418, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N420, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N422, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N424, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N426, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N428, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N430, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N432, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N434, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N436, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N438, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N440, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N442, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N444, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N446, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N448, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N450, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N452, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N454, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N456, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N458, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N460, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N462, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N464, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N466, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N468, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N470, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N472, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N411, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N413, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N415, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N417, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N419, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N421, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N423, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N425, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N427, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N429, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N431, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N433, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N435, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N437, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N439, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N441, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N443, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N445, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N447, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N449, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N451, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N453, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N455, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N457, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N459, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N461, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N463, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N465, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N467, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N469, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N471, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N473, 
         -- Connections to port 'Z'
         Z(0) => N556 );
   C13245_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_13_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_13_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_13_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_13_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_13_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_13_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_13_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_13_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_13_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_13_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_13_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_13_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_13_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_13_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_13_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_13_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_13_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_13_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_13_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_13_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_13_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_13_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_13_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_13_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_13_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_13_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_13_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_13_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_13_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_13_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_13_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_13_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_13_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_13_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_13_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_13_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_13_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_13_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_13_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_13_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_13_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_13_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_13_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_13_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_13_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_13_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_13_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_13_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_13_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_13_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_13_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_13_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_13_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_13_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_13_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_13_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_13_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_13_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_13_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_13_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_13_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_13_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_13_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_13_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N410, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N412, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N414, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N416, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N418, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N420, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N422, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N424, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N426, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N428, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N430, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N432, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N434, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N436, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N438, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N440, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N442, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N444, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N446, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N448, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N450, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N452, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N454, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N456, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N458, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N460, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N462, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N464, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N466, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N468, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N470, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N472, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N411, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N413, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N415, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N417, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N419, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N421, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N423, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N425, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N427, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N429, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N431, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N433, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N435, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N437, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N439, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N441, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N443, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N445, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N447, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N449, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N451, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N453, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N455, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N457, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N459, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N461, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N463, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N465, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N467, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N469, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N471, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N473, 
         -- Connections to port 'Z'
         Z(0) => N557 );
   C13246_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_12_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_12_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_12_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_12_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_12_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_12_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_12_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_12_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_12_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_12_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_12_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_12_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_12_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_12_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_12_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_12_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_12_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_12_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_12_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_12_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_12_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_12_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_12_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_12_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_12_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_12_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_12_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_12_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_12_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_12_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_12_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_12_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_12_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_12_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_12_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_12_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_12_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_12_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_12_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_12_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_12_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_12_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_12_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_12_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_12_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_12_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_12_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_12_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_12_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_12_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_12_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_12_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_12_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_12_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_12_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_12_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_12_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_12_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_12_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_12_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_12_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_12_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_12_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_12_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N410, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N412, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N414, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N416, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N418, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N420, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N422, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N424, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N426, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N428, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N430, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N432, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N434, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N436, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N438, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N440, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N442, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N444, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N446, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N448, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N450, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N452, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N454, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N456, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N458, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N460, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N462, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N464, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N466, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N468, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N470, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N472, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N411, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N413, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N415, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N417, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N419, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N421, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N423, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N425, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N427, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N429, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N431, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N433, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N435, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N437, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N439, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N441, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N443, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N445, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N447, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N449, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N451, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N453, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N455, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N457, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N459, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N461, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N463, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N465, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N467, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N469, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N471, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N473, 
         -- Connections to port 'Z'
         Z(0) => N558 );
   C13247_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_11_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_11_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_11_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_11_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_11_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_11_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_11_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_11_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_11_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_11_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_11_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_11_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_11_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_11_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_11_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_11_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_11_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_11_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_11_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_11_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_11_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_11_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_11_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_11_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_11_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_11_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_11_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_11_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_11_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_11_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_11_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_11_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_11_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_11_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_11_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_11_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_11_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_11_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_11_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_11_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_11_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_11_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_11_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_11_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_11_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_11_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_11_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_11_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_11_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_11_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_11_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_11_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_11_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_11_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_11_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_11_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_11_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_11_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_11_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_11_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_11_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_11_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_11_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_11_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N410, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N412, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N414, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N416, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N418, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N420, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N422, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N424, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N426, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N428, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N430, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N432, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N434, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N436, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N438, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N440, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N442, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N444, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N446, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N448, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N450, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N452, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N454, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N456, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N458, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N460, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N462, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N464, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N466, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N468, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N470, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N472, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N411, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N413, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N415, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N417, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N419, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N421, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N423, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N425, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N427, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N429, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N431, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N433, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N435, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N437, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N439, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N441, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N443, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N445, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N447, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N449, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N451, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N453, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N455, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N457, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N459, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N461, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N463, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N465, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N467, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N469, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N471, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N473, 
         -- Connections to port 'Z'
         Z(0) => N559 );
   C13248_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_10_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_10_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_10_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_10_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_10_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_10_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_10_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_10_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_10_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_10_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_10_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_10_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_10_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_10_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_10_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_10_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_10_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_10_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_10_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_10_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_10_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_10_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_10_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_10_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_10_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_10_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_10_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_10_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_10_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_10_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_10_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_10_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_10_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_10_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_10_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_10_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_10_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_10_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_10_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_10_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_10_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_10_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_10_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_10_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_10_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_10_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_10_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_10_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_10_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_10_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_10_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_10_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_10_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_10_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_10_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_10_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_10_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_10_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_10_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_10_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_10_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_10_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_10_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_10_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N410, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N412, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N414, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N416, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N418, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N420, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N422, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N424, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N426, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N428, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N430, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N432, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N434, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N436, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N438, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N440, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N442, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N444, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N446, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N448, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N450, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N452, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N454, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N456, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N458, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N460, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N462, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N464, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N466, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N468, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N470, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N472, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N411, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N413, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N415, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N417, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N419, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N421, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N423, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N425, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N427, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N429, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N431, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N433, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N435, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N437, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N439, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N441, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N443, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N445, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N447, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N449, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N451, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N453, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N455, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N457, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N459, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N461, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N463, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N465, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N467, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N469, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N471, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N473, 
         -- Connections to port 'Z'
         Z(0) => N560 );
   C13249_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_9_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_9_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_9_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_9_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_9_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_9_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_9_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_9_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_9_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_9_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_9_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_9_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_9_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_9_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_9_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_9_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_9_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_9_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_9_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_9_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_9_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_9_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_9_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_9_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_9_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_9_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_9_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_9_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_9_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_9_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_9_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_9_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_9_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_9_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_9_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_9_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_9_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_9_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_9_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_9_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_9_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_9_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_9_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_9_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_9_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_9_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_9_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_9_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_9_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_9_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_9_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_9_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_9_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_9_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_9_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_9_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_9_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_9_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_9_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_9_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_9_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_9_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_9_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_9_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N410, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N412, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N414, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N416, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N418, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N420, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N422, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N424, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N426, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N428, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N430, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N432, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N434, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N436, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N438, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N440, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N442, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N444, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N446, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N448, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N450, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N452, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N454, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N456, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N458, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N460, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N462, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N464, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N466, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N468, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N470, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N472, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N411, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N413, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N415, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N417, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N419, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N421, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N423, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N425, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N427, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N429, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N431, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N433, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N435, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N437, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N439, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N441, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N443, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N445, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N447, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N449, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N451, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N453, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N455, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N457, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N459, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N461, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N463, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N465, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N467, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N469, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N471, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N473, 
         -- Connections to port 'Z'
         Z(0) => N561 );
   C13250_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_8_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_8_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_8_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_8_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_8_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_8_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_8_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_8_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_8_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_8_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_8_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_8_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_8_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_8_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_8_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_8_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_8_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_8_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_8_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_8_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_8_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_8_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_8_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_8_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_8_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_8_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_8_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_8_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_8_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_8_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_8_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_8_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_8_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_8_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_8_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_8_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_8_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_8_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_8_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_8_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_8_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_8_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_8_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_8_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_8_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_8_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_8_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_8_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_8_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_8_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_8_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_8_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_8_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_8_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_8_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_8_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_8_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_8_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_8_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_8_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_8_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_8_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_8_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_8_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N410, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N412, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N414, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N416, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N418, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N420, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N422, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N424, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N426, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N428, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N430, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N432, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N434, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N436, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N438, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N440, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N442, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N444, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N446, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N448, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N450, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N452, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N454, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N456, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N458, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N460, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N462, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N464, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N466, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N468, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N470, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N472, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N411, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N413, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N415, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N417, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N419, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N421, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N423, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N425, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N427, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N429, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N431, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N433, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N435, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N437, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N439, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N441, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N443, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N445, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N447, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N449, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N451, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N453, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N455, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N457, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N459, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N461, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N463, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N465, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N467, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N469, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N471, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N473, 
         -- Connections to port 'Z'
         Z(0) => N562 );
   C13251_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_7_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_7_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_7_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_7_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_7_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_7_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_7_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_7_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_7_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_7_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_7_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_7_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_7_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_7_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_7_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_7_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_7_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_7_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_7_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_7_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_7_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_7_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_7_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_7_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_7_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_7_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_7_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_7_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_7_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_7_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_7_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_7_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_7_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_7_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_7_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_7_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_7_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_7_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_7_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_7_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_7_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_7_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_7_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_7_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_7_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_7_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_7_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_7_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_7_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_7_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_7_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_7_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_7_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_7_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_7_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_7_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_7_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_7_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_7_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_7_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_7_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_7_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_7_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_7_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N410, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N412, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N414, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N416, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N418, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N420, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N422, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N424, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N426, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N428, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N430, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N432, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N434, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N436, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N438, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N440, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N442, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N444, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N446, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N448, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N450, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N452, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N454, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N456, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N458, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N460, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N462, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N464, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N466, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N468, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N470, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N472, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N411, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N413, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N415, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N417, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N419, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N421, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N423, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N425, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N427, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N429, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N431, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N433, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N435, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N437, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N439, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N441, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N443, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N445, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N447, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N449, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N451, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N453, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N455, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N457, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N459, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N461, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N463, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N465, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N467, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N469, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N471, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N473, 
         -- Connections to port 'Z'
         Z(0) => N563 );
   C13252_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_6_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_6_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_6_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_6_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_6_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_6_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_6_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_6_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_6_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_6_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_6_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_6_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_6_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_6_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_6_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_6_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_6_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_6_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_6_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_6_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_6_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_6_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_6_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_6_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_6_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_6_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_6_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_6_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_6_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_6_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_6_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_6_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_6_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_6_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_6_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_6_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_6_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_6_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_6_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_6_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_6_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_6_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_6_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_6_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_6_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_6_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_6_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_6_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_6_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_6_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_6_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_6_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_6_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_6_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_6_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_6_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_6_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_6_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_6_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_6_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_6_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_6_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_6_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_6_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N410, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N412, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N414, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N416, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N418, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N420, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N422, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N424, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N426, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N428, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N430, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N432, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N434, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N436, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N438, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N440, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N442, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N444, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N446, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N448, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N450, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N452, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N454, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N456, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N458, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N460, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N462, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N464, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N466, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N468, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N470, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N472, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N411, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N413, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N415, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N417, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N419, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N421, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N423, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N425, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N427, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N429, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N431, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N433, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N435, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N437, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N439, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N441, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N443, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N445, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N447, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N449, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N451, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N453, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N455, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N457, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N459, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N461, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N463, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N465, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N467, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N469, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N471, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N473, 
         -- Connections to port 'Z'
         Z(0) => N564 );
   C13253_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_5_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_5_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_5_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_5_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_5_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_5_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_5_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_5_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_5_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_5_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_5_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_5_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_5_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_5_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_5_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_5_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_5_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_5_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_5_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_5_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_5_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_5_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_5_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_5_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_5_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_5_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_5_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_5_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_5_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_5_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_5_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_5_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_5_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_5_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_5_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_5_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_5_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_5_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_5_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_5_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_5_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_5_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_5_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_5_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_5_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_5_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_5_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_5_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_5_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_5_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_5_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_5_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_5_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_5_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_5_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_5_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_5_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_5_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_5_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_5_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_5_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_5_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_5_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_5_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N410, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N412, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N414, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N416, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N418, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N420, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N422, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N424, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N426, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N428, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N430, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N432, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N434, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N436, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N438, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N440, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N442, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N444, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N446, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N448, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N450, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N452, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N454, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N456, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N458, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N460, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N462, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N464, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N466, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N468, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N470, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N472, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N411, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N413, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N415, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N417, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N419, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N421, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N423, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N425, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N427, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N429, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N431, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N433, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N435, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N437, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N439, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N441, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N443, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N445, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N447, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N449, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N451, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N453, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N455, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N457, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N459, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N461, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N463, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N465, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N467, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N469, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N471, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N473, 
         -- Connections to port 'Z'
         Z(0) => N565 );
   C13254_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_4_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_4_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_4_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_4_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_4_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_4_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_4_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_4_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_4_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_4_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_4_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_4_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_4_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_4_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_4_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_4_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_4_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_4_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_4_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_4_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_4_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_4_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_4_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_4_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_4_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_4_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_4_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_4_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_4_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_4_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_4_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_4_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_4_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_4_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_4_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_4_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_4_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_4_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_4_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_4_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_4_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_4_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_4_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_4_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_4_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_4_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_4_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_4_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_4_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_4_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_4_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_4_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_4_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_4_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_4_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_4_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_4_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_4_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_4_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_4_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_4_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_4_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_4_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_4_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N410, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N412, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N414, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N416, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N418, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N420, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N422, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N424, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N426, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N428, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N430, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N432, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N434, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N436, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N438, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N440, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N442, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N444, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N446, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N448, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N450, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N452, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N454, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N456, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N458, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N460, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N462, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N464, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N466, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N468, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N470, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N472, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N411, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N413, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N415, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N417, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N419, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N421, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N423, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N425, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N427, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N429, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N431, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N433, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N435, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N437, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N439, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N441, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N443, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N445, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N447, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N449, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N451, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N453, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N455, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N457, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N459, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N461, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N463, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N465, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N467, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N469, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N471, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N473, 
         -- Connections to port 'Z'
         Z(0) => N566 );
   C13255_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_3_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_3_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_3_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_3_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_3_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_3_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_3_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_3_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_3_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_3_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_3_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_3_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_3_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_3_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_3_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_3_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_3_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_3_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_3_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_3_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_3_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_3_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_3_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_3_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_3_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_3_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_3_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_3_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_3_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_3_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_3_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_3_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_3_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_3_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_3_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_3_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_3_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_3_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_3_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_3_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_3_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_3_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_3_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_3_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_3_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_3_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_3_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_3_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_3_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_3_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_3_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_3_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_3_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_3_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_3_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_3_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_3_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_3_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_3_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_3_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_3_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_3_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_3_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_3_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N410, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N412, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N414, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N416, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N418, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N420, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N422, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N424, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N426, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N428, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N430, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N432, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N434, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N436, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N438, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N440, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N442, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N444, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N446, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N448, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N450, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N452, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N454, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N456, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N458, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N460, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N462, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N464, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N466, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N468, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N470, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N472, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N411, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N413, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N415, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N417, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N419, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N421, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N423, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N425, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N427, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N429, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N431, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N433, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N435, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N437, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N439, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N441, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N443, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N445, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N447, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N449, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N451, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N453, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N455, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N457, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N459, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N461, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N463, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N465, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N467, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N469, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N471, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N473, 
         -- Connections to port 'Z'
         Z(0) => N567 );
   C13256_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_2_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_2_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_2_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_2_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_2_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_2_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_2_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_2_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_2_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_2_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_2_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_2_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_2_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_2_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_2_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_2_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_2_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_2_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_2_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_2_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_2_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_2_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_2_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_2_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_2_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_2_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_2_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_2_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_2_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_2_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_2_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_2_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_2_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_2_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_2_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_2_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_2_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_2_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_2_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_2_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_2_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_2_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_2_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_2_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_2_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_2_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_2_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_2_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_2_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_2_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_2_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_2_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_2_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_2_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_2_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_2_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_2_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_2_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_2_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_2_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_2_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_2_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_2_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_2_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N410, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N412, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N414, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N416, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N418, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N420, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N422, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N424, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N426, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N428, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N430, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N432, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N434, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N436, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N438, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N440, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N442, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N444, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N446, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N448, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N450, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N452, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N454, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N456, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N458, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N460, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N462, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N464, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N466, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N468, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N470, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N472, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N411, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N413, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N415, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N417, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N419, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N421, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N423, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N425, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N427, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N429, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N431, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N433, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N435, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N437, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N439, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N441, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N443, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N445, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N447, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N449, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N451, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N453, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N455, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N457, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N459, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N461, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N463, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N465, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N467, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N469, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N471, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N473, 
         -- Connections to port 'Z'
         Z(0) => N568 );
   C13257_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_1_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_1_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_1_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_1_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_1_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_1_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_1_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_1_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_1_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_1_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_1_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_1_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_1_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_1_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_1_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_1_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_1_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_1_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_1_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_1_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_1_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_1_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_1_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_1_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_1_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_1_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_1_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_1_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_1_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_1_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_1_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_1_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_1_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_1_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_1_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_1_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_1_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_1_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_1_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_1_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_1_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_1_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_1_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_1_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_1_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_1_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_1_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_1_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_1_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_1_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_1_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_1_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_1_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_1_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_1_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_1_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_1_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_1_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_1_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_1_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_1_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_1_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_1_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_1_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N410, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N412, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N414, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N416, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N418, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N420, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N422, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N424, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N426, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N428, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N430, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N432, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N434, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N436, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N438, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N440, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N442, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N444, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N446, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N448, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N450, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N452, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N454, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N456, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N458, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N460, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N462, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N464, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N466, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N468, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N470, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N472, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N411, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N413, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N415, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N417, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N419, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N421, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N423, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N425, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N427, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N429, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N431, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N433, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N435, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N437, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N439, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N441, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N443, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N445, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N447, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N449, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N451, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N453, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N455, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N457, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N459, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N461, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N463, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N465, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N467, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N469, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N471, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N473, 
         -- Connections to port 'Z'
         Z(0) => N569 );
   C13258_cell : SELECT_OP
      generic map ( num_inputs => 64, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_0_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_0_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_0_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_0_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_0_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_0_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_0_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_0_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_0_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_0_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_0_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_0_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_0_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_0_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_0_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_0_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_0_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_0_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_0_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_0_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_0_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_0_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_0_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_0_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_0_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_0_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_0_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_0_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_0_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_0_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_0_port, 
         -- Connections to port 'DATA33'
         DATA(32) => REGISTERS_32_0_port, 
         -- Connections to port 'DATA34'
         DATA(33) => REGISTERS_33_0_port, 
         -- Connections to port 'DATA35'
         DATA(34) => REGISTERS_34_0_port, 
         -- Connections to port 'DATA36'
         DATA(35) => REGISTERS_35_0_port, 
         -- Connections to port 'DATA37'
         DATA(36) => REGISTERS_36_0_port, 
         -- Connections to port 'DATA38'
         DATA(37) => REGISTERS_37_0_port, 
         -- Connections to port 'DATA39'
         DATA(38) => REGISTERS_38_0_port, 
         -- Connections to port 'DATA40'
         DATA(39) => REGISTERS_39_0_port, 
         -- Connections to port 'DATA41'
         DATA(40) => REGISTERS_40_0_port, 
         -- Connections to port 'DATA42'
         DATA(41) => REGISTERS_41_0_port, 
         -- Connections to port 'DATA43'
         DATA(42) => REGISTERS_42_0_port, 
         -- Connections to port 'DATA44'
         DATA(43) => REGISTERS_43_0_port, 
         -- Connections to port 'DATA45'
         DATA(44) => REGISTERS_44_0_port, 
         -- Connections to port 'DATA46'
         DATA(45) => REGISTERS_45_0_port, 
         -- Connections to port 'DATA47'
         DATA(46) => REGISTERS_46_0_port, 
         -- Connections to port 'DATA48'
         DATA(47) => REGISTERS_47_0_port, 
         -- Connections to port 'DATA49'
         DATA(48) => REGISTERS_48_0_port, 
         -- Connections to port 'DATA50'
         DATA(49) => REGISTERS_49_0_port, 
         -- Connections to port 'DATA51'
         DATA(50) => REGISTERS_50_0_port, 
         -- Connections to port 'DATA52'
         DATA(51) => REGISTERS_51_0_port, 
         -- Connections to port 'DATA53'
         DATA(52) => REGISTERS_52_0_port, 
         -- Connections to port 'DATA54'
         DATA(53) => REGISTERS_53_0_port, 
         -- Connections to port 'DATA55'
         DATA(54) => REGISTERS_54_0_port, 
         -- Connections to port 'DATA56'
         DATA(55) => REGISTERS_55_0_port, 
         -- Connections to port 'DATA57'
         DATA(56) => REGISTERS_56_0_port, 
         -- Connections to port 'DATA58'
         DATA(57) => REGISTERS_57_0_port, 
         -- Connections to port 'DATA59'
         DATA(58) => REGISTERS_58_0_port, 
         -- Connections to port 'DATA60'
         DATA(59) => REGISTERS_59_0_port, 
         -- Connections to port 'DATA61'
         DATA(60) => REGISTERS_60_0_port, 
         -- Connections to port 'DATA62'
         DATA(61) => REGISTERS_61_0_port, 
         -- Connections to port 'DATA63'
         DATA(62) => REGISTERS_62_0_port, 
         -- Connections to port 'DATA64'
         DATA(63) => REGISTERS_63_0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N410, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N412, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N414, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N416, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N418, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N420, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N422, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N424, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N426, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N428, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N430, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N432, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N434, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N436, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N438, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N440, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N442, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N444, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N446, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N448, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N450, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N452, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N454, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N456, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N458, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N460, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N462, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N464, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N466, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N468, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N470, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N472, 
         -- Connections to port 'CONTROL33'
         CONTROL(32) => N411, 
         -- Connections to port 'CONTROL34'
         CONTROL(33) => N413, 
         -- Connections to port 'CONTROL35'
         CONTROL(34) => N415, 
         -- Connections to port 'CONTROL36'
         CONTROL(35) => N417, 
         -- Connections to port 'CONTROL37'
         CONTROL(36) => N419, 
         -- Connections to port 'CONTROL38'
         CONTROL(37) => N421, 
         -- Connections to port 'CONTROL39'
         CONTROL(38) => N423, 
         -- Connections to port 'CONTROL40'
         CONTROL(39) => N425, 
         -- Connections to port 'CONTROL41'
         CONTROL(40) => N427, 
         -- Connections to port 'CONTROL42'
         CONTROL(41) => N429, 
         -- Connections to port 'CONTROL43'
         CONTROL(42) => N431, 
         -- Connections to port 'CONTROL44'
         CONTROL(43) => N433, 
         -- Connections to port 'CONTROL45'
         CONTROL(44) => N435, 
         -- Connections to port 'CONTROL46'
         CONTROL(45) => N437, 
         -- Connections to port 'CONTROL47'
         CONTROL(46) => N439, 
         -- Connections to port 'CONTROL48'
         CONTROL(47) => N441, 
         -- Connections to port 'CONTROL49'
         CONTROL(48) => N443, 
         -- Connections to port 'CONTROL50'
         CONTROL(49) => N445, 
         -- Connections to port 'CONTROL51'
         CONTROL(50) => N447, 
         -- Connections to port 'CONTROL52'
         CONTROL(51) => N449, 
         -- Connections to port 'CONTROL53'
         CONTROL(52) => N451, 
         -- Connections to port 'CONTROL54'
         CONTROL(53) => N453, 
         -- Connections to port 'CONTROL55'
         CONTROL(54) => N455, 
         -- Connections to port 'CONTROL56'
         CONTROL(55) => N457, 
         -- Connections to port 'CONTROL57'
         CONTROL(56) => N459, 
         -- Connections to port 'CONTROL58'
         CONTROL(57) => N461, 
         -- Connections to port 'CONTROL59'
         CONTROL(58) => N463, 
         -- Connections to port 'CONTROL60'
         CONTROL(59) => N465, 
         -- Connections to port 'CONTROL61'
         CONTROL(60) => N467, 
         -- Connections to port 'CONTROL62'
         CONTROL(61) => N469, 
         -- Connections to port 'CONTROL63'
         CONTROL(62) => N471, 
         -- Connections to port 'CONTROL64'
         CONTROL(63) => N473, 
         -- Connections to port 'Z'
         Z(0) => N570 );
   OUT1_reg_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N638, next_state => N604, 
               clocked_on => CLK_port, Q => OUT1_31_port, QN => n_3048);
   OUT1_reg_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N638, next_state => N603, 
               clocked_on => CLK_port, Q => OUT1_30_port, QN => n_3049);
   OUT1_reg_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N638, next_state => N602, 
               clocked_on => CLK_port, Q => OUT1_29_port, QN => n_3050);
   OUT1_reg_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N638, next_state => N601, 
               clocked_on => CLK_port, Q => OUT1_28_port, QN => n_3051);
   OUT1_reg_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N638, next_state => N600, 
               clocked_on => CLK_port, Q => OUT1_27_port, QN => n_3052);
   OUT1_reg_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N638, next_state => N599, 
               clocked_on => CLK_port, Q => OUT1_26_port, QN => n_3053);
   OUT1_reg_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N638, next_state => N598, 
               clocked_on => CLK_port, Q => OUT1_25_port, QN => n_3054);
   OUT1_reg_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N638, next_state => N597, 
               clocked_on => CLK_port, Q => OUT1_24_port, QN => n_3055);
   OUT1_reg_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N638, next_state => N596, 
               clocked_on => CLK_port, Q => OUT1_23_port, QN => n_3056);
   OUT1_reg_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N638, next_state => N595, 
               clocked_on => CLK_port, Q => OUT1_22_port, QN => n_3057);
   OUT1_reg_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N638, next_state => N594, 
               clocked_on => CLK_port, Q => OUT1_21_port, QN => n_3058);
   OUT1_reg_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N638, next_state => N593, 
               clocked_on => CLK_port, Q => OUT1_20_port, QN => n_3059);
   OUT1_reg_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N638, next_state => N592, 
               clocked_on => CLK_port, Q => OUT1_19_port, QN => n_3060);
   OUT1_reg_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N638, next_state => N591, 
               clocked_on => CLK_port, Q => OUT1_18_port, QN => n_3061);
   OUT1_reg_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N638, next_state => N590, 
               clocked_on => CLK_port, Q => OUT1_17_port, QN => n_3062);
   OUT1_reg_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N638, next_state => N589, 
               clocked_on => CLK_port, Q => OUT1_16_port, QN => n_3063);
   OUT1_reg_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N638, next_state => N588, 
               clocked_on => CLK_port, Q => OUT1_15_port, QN => n_3064);
   OUT1_reg_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N638, next_state => N587, 
               clocked_on => CLK_port, Q => OUT1_14_port, QN => n_3065);
   OUT1_reg_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N638, next_state => N586, 
               clocked_on => CLK_port, Q => OUT1_13_port, QN => n_3066);
   OUT1_reg_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N638, next_state => N585, 
               clocked_on => CLK_port, Q => OUT1_12_port, QN => n_3067);
   OUT1_reg_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N638, next_state => N584, 
               clocked_on => CLK_port, Q => OUT1_11_port, QN => n_3068);
   OUT1_reg_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N638, next_state => N583, 
               clocked_on => CLK_port, Q => OUT1_10_port, QN => n_3069);
   OUT1_reg_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N638, next_state => N582, 
               clocked_on => CLK_port, Q => OUT1_9_port, QN => n_3070);
   OUT1_reg_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N638, next_state => N581, 
               clocked_on => CLK_port, Q => OUT1_8_port, QN => n_3071);
   OUT1_reg_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N638, next_state => N580, 
               clocked_on => CLK_port, Q => OUT1_7_port, QN => n_3072);
   OUT1_reg_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N638, next_state => N579, 
               clocked_on => CLK_port, Q => OUT1_6_port, QN => n_3073);
   OUT1_reg_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N638, next_state => N578, 
               clocked_on => CLK_port, Q => OUT1_5_port, QN => n_3074);
   OUT1_reg_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N638, next_state => N577, 
               clocked_on => CLK_port, Q => OUT1_4_port, QN => n_3075);
   OUT1_reg_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N638, next_state => N576, 
               clocked_on => CLK_port, Q => OUT1_3_port, QN => n_3076);
   OUT1_reg_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N638, next_state => N575, 
               clocked_on => CLK_port, Q => OUT1_2_port, QN => n_3077);
   OUT1_reg_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N638, next_state => N574, 
               clocked_on => CLK_port, Q => OUT1_1_port, QN => n_3078);
   OUT1_reg_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N638, next_state => N573, 
               clocked_on => CLK_port, Q => OUT1_0_port, QN => n_3079);
   OUT2_reg_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N639, next_state => N637, 
               clocked_on => CLK_port, Q => OUT2_31_port, QN => n_3080);
   OUT2_reg_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N639, next_state => N636, 
               clocked_on => CLK_port, Q => OUT2_30_port, QN => n_3081);
   OUT2_reg_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N639, next_state => N635, 
               clocked_on => CLK_port, Q => OUT2_29_port, QN => n_3082);
   OUT2_reg_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N639, next_state => N634, 
               clocked_on => CLK_port, Q => OUT2_28_port, QN => n_3083);
   OUT2_reg_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N639, next_state => N633, 
               clocked_on => CLK_port, Q => OUT2_27_port, QN => n_3084);
   OUT2_reg_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N639, next_state => N632, 
               clocked_on => CLK_port, Q => OUT2_26_port, QN => n_3085);
   OUT2_reg_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N639, next_state => N631, 
               clocked_on => CLK_port, Q => OUT2_25_port, QN => n_3086);
   OUT2_reg_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N639, next_state => N630, 
               clocked_on => CLK_port, Q => OUT2_24_port, QN => n_3087);
   OUT2_reg_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N639, next_state => N629, 
               clocked_on => CLK_port, Q => OUT2_23_port, QN => n_3088);
   OUT2_reg_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N639, next_state => N628, 
               clocked_on => CLK_port, Q => OUT2_22_port, QN => n_3089);
   OUT2_reg_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N639, next_state => N627, 
               clocked_on => CLK_port, Q => OUT2_21_port, QN => n_3090);
   OUT2_reg_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N639, next_state => N626, 
               clocked_on => CLK_port, Q => OUT2_20_port, QN => n_3091);
   OUT2_reg_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N639, next_state => N625, 
               clocked_on => CLK_port, Q => OUT2_19_port, QN => n_3092);
   OUT2_reg_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N639, next_state => N624, 
               clocked_on => CLK_port, Q => OUT2_18_port, QN => n_3093);
   OUT2_reg_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N639, next_state => N623, 
               clocked_on => CLK_port, Q => OUT2_17_port, QN => n_3094);
   OUT2_reg_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N639, next_state => N622, 
               clocked_on => CLK_port, Q => OUT2_16_port, QN => n_3095);
   OUT2_reg_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N639, next_state => N621, 
               clocked_on => CLK_port, Q => OUT2_15_port, QN => n_3096);
   OUT2_reg_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N639, next_state => N620, 
               clocked_on => CLK_port, Q => OUT2_14_port, QN => n_3097);
   OUT2_reg_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N639, next_state => N619, 
               clocked_on => CLK_port, Q => OUT2_13_port, QN => n_3098);
   OUT2_reg_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N639, next_state => N618, 
               clocked_on => CLK_port, Q => OUT2_12_port, QN => n_3099);
   OUT2_reg_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N639, next_state => N617, 
               clocked_on => CLK_port, Q => OUT2_11_port, QN => n_3100);
   OUT2_reg_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N639, next_state => N616, 
               clocked_on => CLK_port, Q => OUT2_10_port, QN => n_3101);
   OUT2_reg_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N639, next_state => N615, 
               clocked_on => CLK_port, Q => OUT2_9_port, QN => n_3102);
   OUT2_reg_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N639, next_state => N614, 
               clocked_on => CLK_port, Q => OUT2_8_port, QN => n_3103);
   OUT2_reg_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N639, next_state => N613, 
               clocked_on => CLK_port, Q => OUT2_7_port, QN => n_3104);
   OUT2_reg_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N639, next_state => N612, 
               clocked_on => CLK_port, Q => OUT2_6_port, QN => n_3105);
   OUT2_reg_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N639, next_state => N611, 
               clocked_on => CLK_port, Q => OUT2_5_port, QN => n_3106);
   OUT2_reg_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N639, next_state => N610, 
               clocked_on => CLK_port, Q => OUT2_4_port, QN => n_3107);
   OUT2_reg_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N639, next_state => N609, 
               clocked_on => CLK_port, Q => OUT2_3_port, QN => n_3108);
   OUT2_reg_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N639, next_state => N608, 
               clocked_on => CLK_port, Q => OUT2_2_port, QN => n_3109);
   OUT2_reg_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N639, next_state => N607, 
               clocked_on => CLK_port, Q => OUT2_1_port, QN => n_3110);
   OUT2_reg_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N639, next_state => N606, 
               clocked_on => CLK_port, Q => OUT2_0_port, QN => n_3111);
   I_0 : GTECH_NOT port map( A => ADD_WR(5), Z => N640);
   C13843 : GTECH_AND2 port map( A => ADD_WR(3), B => ADD_WR(4), Z => N641);
   C13844 : GTECH_AND2 port map( A => N0, B => ADD_WR(4), Z => N642);
   I_1 : GTECH_NOT port map( A => ADD_WR(3), Z => N0);
   C13845 : GTECH_AND2 port map( A => ADD_WR(3), B => N1, Z => N643);
   I_2 : GTECH_NOT port map( A => ADD_WR(4), Z => N1);
   C13846 : GTECH_AND2 port map( A => N2, B => N3, Z => N644);
   I_3 : GTECH_NOT port map( A => ADD_WR(3), Z => N2);
   I_4 : GTECH_NOT port map( A => ADD_WR(4), Z => N3);
   C13847 : GTECH_AND2 port map( A => ADD_WR(5), B => N641, Z => N645);
   C13848 : GTECH_AND2 port map( A => ADD_WR(5), B => N642, Z => N646);
   C13849 : GTECH_AND2 port map( A => ADD_WR(5), B => N643, Z => N647);
   C13850 : GTECH_AND2 port map( A => ADD_WR(5), B => N644, Z => N648);
   C13851 : GTECH_AND2 port map( A => N640, B => N641, Z => N649);
   C13852 : GTECH_AND2 port map( A => N640, B => N642, Z => N650);
   C13853 : GTECH_AND2 port map( A => N640, B => N643, Z => N651);
   C13854 : GTECH_AND2 port map( A => N640, B => N644, Z => N652);
   I_5 : GTECH_NOT port map( A => ADD_WR(2), Z => N653);
   C13856 : GTECH_AND2 port map( A => ADD_WR(0), B => ADD_WR(1), Z => N654);
   C13857 : GTECH_AND2 port map( A => N4, B => ADD_WR(1), Z => N655);
   I_6 : GTECH_NOT port map( A => ADD_WR(0), Z => N4);
   C13858 : GTECH_AND2 port map( A => ADD_WR(0), B => N5, Z => N656);
   I_7 : GTECH_NOT port map( A => ADD_WR(1), Z => N5);
   C13859 : GTECH_AND2 port map( A => N6, B => N7, Z => N657);
   I_8 : GTECH_NOT port map( A => ADD_WR(0), Z => N6);
   I_9 : GTECH_NOT port map( A => ADD_WR(1), Z => N7);
   C13860 : GTECH_AND2 port map( A => ADD_WR(2), B => N654, Z => N658);
   C13861 : GTECH_AND2 port map( A => ADD_WR(2), B => N655, Z => N659);
   C13862 : GTECH_AND2 port map( A => ADD_WR(2), B => N656, Z => N660);
   C13863 : GTECH_AND2 port map( A => ADD_WR(2), B => N657, Z => N661);
   C13864 : GTECH_AND2 port map( A => N653, B => N654, Z => N662);
   C13865 : GTECH_AND2 port map( A => N653, B => N655, Z => N663);
   C13866 : GTECH_AND2 port map( A => N653, B => N656, Z => N664);
   C13867 : GTECH_AND2 port map( A => N653, B => N657, Z => N665);
   C13868 : GTECH_AND2 port map( A => N645, B => N658, Z => N666);
   C13869 : GTECH_AND2 port map( A => N645, B => N659, Z => N667);
   C13870 : GTECH_AND2 port map( A => N645, B => N660, Z => N668);
   C13871 : GTECH_AND2 port map( A => N645, B => N661, Z => N669);
   C13872 : GTECH_AND2 port map( A => N645, B => N662, Z => N670);
   C13873 : GTECH_AND2 port map( A => N645, B => N663, Z => N671);
   C13874 : GTECH_AND2 port map( A => N645, B => N664, Z => N672);
   C13875 : GTECH_AND2 port map( A => N645, B => N665, Z => N673);
   C13876 : GTECH_AND2 port map( A => N646, B => N658, Z => N674);
   C13877 : GTECH_AND2 port map( A => N646, B => N659, Z => N675);
   C13878 : GTECH_AND2 port map( A => N646, B => N660, Z => N676);
   C13879 : GTECH_AND2 port map( A => N646, B => N661, Z => N677);
   C13880 : GTECH_AND2 port map( A => N646, B => N662, Z => N678);
   C13881 : GTECH_AND2 port map( A => N646, B => N663, Z => N679);
   C13882 : GTECH_AND2 port map( A => N646, B => N664, Z => N680);
   C13883 : GTECH_AND2 port map( A => N646, B => N665, Z => N681);
   C13884 : GTECH_AND2 port map( A => N647, B => N658, Z => N682);
   C13885 : GTECH_AND2 port map( A => N647, B => N659, Z => N683);
   C13886 : GTECH_AND2 port map( A => N647, B => N660, Z => N684);
   C13887 : GTECH_AND2 port map( A => N647, B => N661, Z => N685);
   C13888 : GTECH_AND2 port map( A => N647, B => N662, Z => N686);
   C13889 : GTECH_AND2 port map( A => N647, B => N663, Z => N687);
   C13890 : GTECH_AND2 port map( A => N647, B => N664, Z => N688);
   C13891 : GTECH_AND2 port map( A => N647, B => N665, Z => N689);
   C13892 : GTECH_AND2 port map( A => N648, B => N658, Z => N690);
   C13893 : GTECH_AND2 port map( A => N648, B => N659, Z => N691);
   C13894 : GTECH_AND2 port map( A => N648, B => N660, Z => N692);
   C13895 : GTECH_AND2 port map( A => N648, B => N661, Z => N693);
   C13896 : GTECH_AND2 port map( A => N648, B => N662, Z => N694);
   C13897 : GTECH_AND2 port map( A => N648, B => N663, Z => N695);
   C13898 : GTECH_AND2 port map( A => N648, B => N664, Z => N696);
   C13899 : GTECH_AND2 port map( A => N648, B => N665, Z => N697);
   C13900 : GTECH_AND2 port map( A => N649, B => N658, Z => N698);
   C13901 : GTECH_AND2 port map( A => N649, B => N659, Z => N699);
   C13902 : GTECH_AND2 port map( A => N649, B => N660, Z => N700);
   C13903 : GTECH_AND2 port map( A => N649, B => N661, Z => N701);
   C13904 : GTECH_AND2 port map( A => N649, B => N662, Z => N702);
   C13905 : GTECH_AND2 port map( A => N649, B => N663, Z => N703);
   C13906 : GTECH_AND2 port map( A => N649, B => N664, Z => N704);
   C13907 : GTECH_AND2 port map( A => N649, B => N665, Z => N705);
   C13908 : GTECH_AND2 port map( A => N650, B => N658, Z => N706);
   C13909 : GTECH_AND2 port map( A => N650, B => N659, Z => N707);
   C13910 : GTECH_AND2 port map( A => N650, B => N660, Z => N708);
   C13911 : GTECH_AND2 port map( A => N650, B => N661, Z => N709);
   C13912 : GTECH_AND2 port map( A => N650, B => N662, Z => N710);
   C13913 : GTECH_AND2 port map( A => N650, B => N663, Z => N711);
   C13914 : GTECH_AND2 port map( A => N650, B => N664, Z => N712);
   C13915 : GTECH_AND2 port map( A => N650, B => N665, Z => N713);
   C13916 : GTECH_AND2 port map( A => N651, B => N658, Z => N714);
   C13917 : GTECH_AND2 port map( A => N651, B => N659, Z => N715);
   C13918 : GTECH_AND2 port map( A => N651, B => N660, Z => N716);
   C13919 : GTECH_AND2 port map( A => N651, B => N661, Z => N717);
   C13920 : GTECH_AND2 port map( A => N651, B => N662, Z => N718);
   C13921 : GTECH_AND2 port map( A => N651, B => N663, Z => N719);
   C13922 : GTECH_AND2 port map( A => N651, B => N664, Z => N720);
   C13923 : GTECH_AND2 port map( A => N651, B => N665, Z => N721);
   C13924 : GTECH_AND2 port map( A => N652, B => N658, Z => N722);
   C13925 : GTECH_AND2 port map( A => N652, B => N659, Z => N723);
   C13926 : GTECH_AND2 port map( A => N652, B => N660, Z => N724);
   C13927 : GTECH_AND2 port map( A => N652, B => N661, Z => N725);
   C13928 : GTECH_AND2 port map( A => N652, B => N662, Z => N726);
   C13929 : GTECH_AND2 port map( A => N652, B => N663, Z => N727);
   C13930 : GTECH_AND2 port map( A => N652, B => N664, Z => N728);
   C13931 : GTECH_AND2 port map( A => N652, B => N665, Z => N729);
   C13932_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 64 )
      port map(
         -- Connections to port 'DATA1'
         DATA(63) => N729, DATA(62) => N728, DATA(61) => N727, DATA(60) => N726
               , DATA(59) => N725, DATA(58) => N724, DATA(57) => N723, DATA(56)
               => N722, DATA(55) => N721, DATA(54) => N720, DATA(53) => N719, 
               DATA(52) => N718, DATA(51) => N717, DATA(50) => N716, DATA(49) 
               => N715, DATA(48) => N714, DATA(47) => N713, DATA(46) => N712, 
               DATA(45) => N711, DATA(44) => N710, DATA(43) => N709, DATA(42) 
               => N708, DATA(41) => N707, DATA(40) => N706, DATA(39) => N705, 
               DATA(38) => N704, DATA(37) => N703, DATA(36) => N702, DATA(35) 
               => N701, DATA(34) => N700, DATA(33) => N699, DATA(32) => N698, 
               DATA(31) => N697, DATA(30) => N696, DATA(29) => N695, DATA(28) 
               => N694, DATA(27) => N693, DATA(26) => N692, DATA(25) => N691, 
               DATA(24) => N690, DATA(23) => N689, DATA(22) => N688, DATA(21) 
               => N687, DATA(20) => N686, DATA(19) => N685, DATA(18) => N684, 
               DATA(17) => N683, DATA(16) => N682, DATA(15) => N681, DATA(14) 
               => N680, DATA(13) => N679, DATA(12) => N678, DATA(11) => N677, 
               DATA(10) => N676, DATA(9) => N675, DATA(8) => N674, DATA(7) => 
               N673, DATA(6) => N672, DATA(5) => N671, DATA(4) => N670, DATA(3)
               => N669, DATA(2) => N668, DATA(1) => N667, DATA(0) => N666, 
         -- Connections to port 'DATA2'
         DATA(127) => X_Logic0_port, DATA(126) => X_Logic0_port, DATA(125) => 
               X_Logic0_port, DATA(124) => X_Logic0_port, DATA(123) => 
               X_Logic0_port, DATA(122) => X_Logic0_port, DATA(121) => 
               X_Logic0_port, DATA(120) => X_Logic0_port, DATA(119) => 
               X_Logic0_port, DATA(118) => X_Logic0_port, DATA(117) => 
               X_Logic0_port, DATA(116) => X_Logic0_port, DATA(115) => 
               X_Logic0_port, DATA(114) => X_Logic0_port, DATA(113) => 
               X_Logic0_port, DATA(112) => X_Logic0_port, DATA(111) => 
               X_Logic0_port, DATA(110) => X_Logic0_port, DATA(109) => 
               X_Logic0_port, DATA(108) => X_Logic0_port, DATA(107) => 
               X_Logic0_port, DATA(106) => X_Logic0_port, DATA(105) => 
               X_Logic0_port, DATA(104) => X_Logic0_port, DATA(103) => 
               X_Logic0_port, DATA(102) => X_Logic0_port, DATA(101) => 
               X_Logic0_port, DATA(100) => X_Logic0_port, DATA(99) => 
               X_Logic0_port, DATA(98) => X_Logic0_port, DATA(97) => 
               X_Logic0_port, DATA(96) => X_Logic0_port, DATA(95) => 
               X_Logic0_port, DATA(94) => X_Logic0_port, DATA(93) => 
               X_Logic0_port, DATA(92) => X_Logic0_port, DATA(91) => 
               X_Logic0_port, DATA(90) => X_Logic0_port, DATA(89) => 
               X_Logic0_port, DATA(88) => X_Logic0_port, DATA(87) => 
               X_Logic0_port, DATA(86) => X_Logic0_port, DATA(85) => 
               X_Logic0_port, DATA(84) => X_Logic0_port, DATA(83) => 
               X_Logic0_port, DATA(82) => X_Logic0_port, DATA(81) => 
               X_Logic0_port, DATA(80) => X_Logic0_port, DATA(79) => 
               X_Logic0_port, DATA(78) => X_Logic0_port, DATA(77) => 
               X_Logic0_port, DATA(76) => X_Logic0_port, DATA(75) => 
               X_Logic0_port, DATA(74) => X_Logic0_port, DATA(73) => 
               X_Logic0_port, DATA(72) => X_Logic0_port, DATA(71) => 
               X_Logic0_port, DATA(70) => X_Logic0_port, DATA(69) => 
               X_Logic0_port, DATA(68) => X_Logic0_port, DATA(67) => 
               X_Logic0_port, DATA(66) => X_Logic0_port, DATA(65) => 
               X_Logic0_port, DATA(64) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N8, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N18, 
         -- Connections to port 'Z'
         Z(63) => N82, Z(62) => N81, Z(61) => N80, Z(60) => N79, Z(59) => N78, 
               Z(58) => N77, Z(57) => N76, Z(56) => N75, Z(55) => N74, Z(54) =>
               N73, Z(53) => N72, Z(52) => N71, Z(51) => N70, Z(50) => N69, 
               Z(49) => N68, Z(48) => N67, Z(47) => N66, Z(46) => N65, Z(45) =>
               N64, Z(44) => N63, Z(43) => N62, Z(42) => N61, Z(41) => N60, 
               Z(40) => N59, Z(39) => N58, Z(38) => N57, Z(37) => N56, Z(36) =>
               N55, Z(35) => N54, Z(34) => N53, Z(33) => N52, Z(32) => N51, 
               Z(31) => N50, Z(30) => N49, Z(29) => N48, Z(28) => N47, Z(27) =>
               N46, Z(26) => N45, Z(25) => N44, Z(24) => N43, Z(23) => N42, 
               Z(22) => N41, Z(21) => N40, Z(20) => N39, Z(19) => N38, Z(18) =>
               N37, Z(17) => N36, Z(16) => N35, Z(15) => N34, Z(14) => N33, 
               Z(13) => N32, Z(12) => N31, Z(11) => N30, Z(10) => N29, Z(9) => 
               N28, Z(8) => N27, Z(7) => N26, Z(6) => N25, Z(5) => N24, Z(4) =>
               N23, Z(3) => N22, Z(2) => N21, Z(1) => N20, Z(0) => N19 );
   B_0 : GTECH_BUF port map( A => N17, Z => N8);
   C13933_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 64 )
      port map(
         -- Connections to port 'DATA1'
         DATA(63) => X_Logic1_port, DATA(62) => X_Logic1_port, DATA(61) => 
               X_Logic1_port, DATA(60) => X_Logic1_port, DATA(59) => 
               X_Logic1_port, DATA(58) => X_Logic1_port, DATA(57) => 
               X_Logic1_port, DATA(56) => X_Logic1_port, DATA(55) => 
               X_Logic1_port, DATA(54) => X_Logic1_port, DATA(53) => 
               X_Logic1_port, DATA(52) => X_Logic1_port, DATA(51) => 
               X_Logic1_port, DATA(50) => X_Logic1_port, DATA(49) => 
               X_Logic1_port, DATA(48) => X_Logic1_port, DATA(47) => 
               X_Logic1_port, DATA(46) => X_Logic1_port, DATA(45) => 
               X_Logic1_port, DATA(44) => X_Logic1_port, DATA(43) => 
               X_Logic1_port, DATA(42) => X_Logic1_port, DATA(41) => 
               X_Logic1_port, DATA(40) => X_Logic1_port, DATA(39) => 
               X_Logic1_port, DATA(38) => X_Logic1_port, DATA(37) => 
               X_Logic1_port, DATA(36) => X_Logic1_port, DATA(35) => 
               X_Logic1_port, DATA(34) => X_Logic1_port, DATA(33) => 
               X_Logic1_port, DATA(32) => X_Logic1_port, DATA(31) => 
               X_Logic1_port, DATA(30) => X_Logic1_port, DATA(29) => 
               X_Logic1_port, DATA(28) => X_Logic1_port, DATA(27) => 
               X_Logic1_port, DATA(26) => X_Logic1_port, DATA(25) => 
               X_Logic1_port, DATA(24) => X_Logic1_port, DATA(23) => 
               X_Logic1_port, DATA(22) => X_Logic1_port, DATA(21) => 
               X_Logic1_port, DATA(20) => X_Logic1_port, DATA(19) => 
               X_Logic1_port, DATA(18) => X_Logic1_port, DATA(17) => 
               X_Logic1_port, DATA(16) => X_Logic1_port, DATA(15) => 
               X_Logic1_port, DATA(14) => X_Logic1_port, DATA(13) => 
               X_Logic1_port, DATA(12) => X_Logic1_port, DATA(11) => 
               X_Logic1_port, DATA(10) => X_Logic1_port, DATA(9) => 
               X_Logic1_port, DATA(8) => X_Logic1_port, DATA(7) => 
               X_Logic1_port, DATA(6) => X_Logic1_port, DATA(5) => 
               X_Logic1_port, DATA(4) => X_Logic1_port, DATA(3) => 
               X_Logic1_port, DATA(2) => X_Logic1_port, DATA(1) => 
               X_Logic1_port, DATA(0) => X_Logic1_port, 
         -- Connections to port 'DATA2'
         DATA(127) => N82, DATA(126) => N81, DATA(125) => N80, DATA(124) => N79
               , DATA(123) => N78, DATA(122) => N77, DATA(121) => N76, 
               DATA(120) => N75, DATA(119) => N74, DATA(118) => N73, DATA(117) 
               => N72, DATA(116) => N71, DATA(115) => N70, DATA(114) => N69, 
               DATA(113) => N68, DATA(112) => N67, DATA(111) => N66, DATA(110) 
               => N65, DATA(109) => N64, DATA(108) => N63, DATA(107) => N62, 
               DATA(106) => N61, DATA(105) => N60, DATA(104) => N59, DATA(103) 
               => N58, DATA(102) => N57, DATA(101) => N56, DATA(100) => N55, 
               DATA(99) => N54, DATA(98) => N53, DATA(97) => N52, DATA(96) => 
               N51, DATA(95) => N50, DATA(94) => N49, DATA(93) => N48, DATA(92)
               => N47, DATA(91) => N46, DATA(90) => N45, DATA(89) => N44, 
               DATA(88) => N43, DATA(87) => N42, DATA(86) => N41, DATA(85) => 
               N40, DATA(84) => N39, DATA(83) => N38, DATA(82) => N37, DATA(81)
               => N36, DATA(80) => N35, DATA(79) => N34, DATA(78) => N33, 
               DATA(77) => N32, DATA(76) => N31, DATA(75) => N30, DATA(74) => 
               N29, DATA(73) => N28, DATA(72) => N27, DATA(71) => N26, DATA(70)
               => N25, DATA(69) => N24, DATA(68) => N23, DATA(67) => N22, 
               DATA(66) => N21, DATA(65) => N20, DATA(64) => N19, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N9, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N10, 
         -- Connections to port 'Z'
         Z(63) => N178, Z(62) => N177, Z(61) => N176, Z(60) => N175, Z(59) => 
               N174, Z(58) => N173, Z(57) => N172, Z(56) => N171, Z(55) => N170
               , Z(54) => N169, Z(53) => N168, Z(52) => N167, Z(51) => N166, 
               Z(50) => N165, Z(49) => N164, Z(48) => N163, Z(47) => N162, 
               Z(46) => N161, Z(45) => N160, Z(44) => N159, Z(43) => N158, 
               Z(42) => N157, Z(41) => N156, Z(40) => N155, Z(39) => N154, 
               Z(38) => N153, Z(37) => N152, Z(36) => N151, Z(35) => N150, 
               Z(34) => N149, Z(33) => N148, Z(32) => N147, Z(31) => N146, 
               Z(30) => N145, Z(29) => N144, Z(28) => N143, Z(27) => N142, 
               Z(26) => N141, Z(25) => N140, Z(24) => N139, Z(23) => N138, 
               Z(22) => N137, Z(21) => N136, Z(20) => N135, Z(19) => N134, 
               Z(18) => N133, Z(17) => N132, Z(16) => N131, Z(15) => N130, 
               Z(14) => N129, Z(13) => N128, Z(12) => N127, Z(11) => N126, 
               Z(10) => N125, Z(9) => N124, Z(8) => N123, Z(7) => N122, Z(6) =>
               N121, Z(5) => N120, Z(4) => N119, Z(3) => N118, Z(2) => N117, 
               Z(1) => N116, Z(0) => N83 );
   B_1 : GTECH_BUF port map( A => RESET, Z => N9);
   B_2 : GTECH_BUF port map( A => N16, Z => N10);
   C13934_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 32 )
      port map(
         -- Connections to port 'DATA1'
         DATA(31) => X_Logic0_port, DATA(30) => X_Logic0_port, DATA(29) => 
               X_Logic0_port, DATA(28) => X_Logic0_port, DATA(27) => 
               X_Logic0_port, DATA(26) => X_Logic0_port, DATA(25) => 
               X_Logic0_port, DATA(24) => X_Logic0_port, DATA(23) => 
               X_Logic0_port, DATA(22) => X_Logic0_port, DATA(21) => 
               X_Logic0_port, DATA(20) => X_Logic0_port, DATA(19) => 
               X_Logic0_port, DATA(18) => X_Logic0_port, DATA(17) => 
               X_Logic0_port, DATA(16) => X_Logic0_port, DATA(15) => 
               X_Logic0_port, DATA(14) => X_Logic0_port, DATA(13) => 
               X_Logic0_port, DATA(12) => X_Logic0_port, DATA(11) => 
               X_Logic0_port, DATA(10) => X_Logic0_port, DATA(9) => 
               X_Logic0_port, DATA(8) => X_Logic0_port, DATA(7) => 
               X_Logic0_port, DATA(6) => X_Logic0_port, DATA(5) => 
               X_Logic0_port, DATA(4) => X_Logic0_port, DATA(3) => 
               X_Logic0_port, DATA(2) => X_Logic0_port, DATA(1) => 
               X_Logic0_port, DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(63) => DATAIN_31_port, DATA(62) => DATAIN_30_port, DATA(61) => 
               DATAIN_29_port, DATA(60) => DATAIN_28_port, DATA(59) => 
               DATAIN_27_port, DATA(58) => DATAIN_26_port, DATA(57) => 
               DATAIN_25_port, DATA(56) => DATAIN_24_port, DATA(55) => 
               DATAIN_23_port, DATA(54) => DATAIN_22_port, DATA(53) => 
               DATAIN_21_port, DATA(52) => DATAIN_20_port, DATA(51) => 
               DATAIN_19_port, DATA(50) => DATAIN_18_port, DATA(49) => 
               DATAIN_17_port, DATA(48) => DATAIN_16_port, DATA(47) => 
               DATAIN_15_port, DATA(46) => DATAIN_14_port, DATA(45) => 
               DATAIN_13_port, DATA(44) => DATAIN_12_port, DATA(43) => 
               DATAIN_11_port, DATA(42) => DATAIN_10_port, DATA(41) => 
               DATAIN_9_port, DATA(40) => DATAIN_8_port, DATA(39) => 
               DATAIN_7_port, DATA(38) => DATAIN_6_port, DATA(37) => 
               DATAIN_5_port, DATA(36) => DATAIN_4_port, DATA(35) => 
               DATAIN_3_port, DATA(34) => DATAIN_2_port, DATA(33) => 
               DATAIN_1_port, DATA(32) => DATAIN_0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N9, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N10, 
         -- Connections to port 'Z'
         Z(31) => N115, Z(30) => N114, Z(29) => N113, Z(28) => N112, Z(27) => 
               N111, Z(26) => N110, Z(25) => N109, Z(24) => N108, Z(23) => N107
               , Z(22) => N106, Z(21) => N105, Z(20) => N104, Z(19) => N103, 
               Z(18) => N102, Z(17) => N101, Z(16) => N100, Z(15) => N99, Z(14)
               => N98, Z(13) => N97, Z(12) => N96, Z(11) => N95, Z(10) => N94, 
               Z(9) => N93, Z(8) => N92, Z(7) => N91, Z(6) => N90, Z(5) => N89,
               Z(4) => N88, Z(3) => N87, Z(2) => N86, Z(1) => N85, Z(0) => N84 
               );
   C13935_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => RD2_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N11, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N12, 
         -- Connections to port 'Z'
         Z(0) => N571 );
   B_3 : GTECH_BUF port map( A => RD1_port, Z => N11);
   B_4 : GTECH_BUF port map( A => N506, Z => N12);
   C13936_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic1_port, 
         -- Connections to port 'DATA2'
         DATA(1) => RD1_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N13, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N181, 
         -- Connections to port 'Z'
         Z(0) => N572 );
   B_5 : GTECH_BUF port map( A => N180, Z => N13);
   C13937_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 32 )
      port map(
         -- Connections to port 'DATA1'
         DATA(31) => N312, DATA(30) => N313, DATA(29) => N314, DATA(28) => N315
               , DATA(27) => N316, DATA(26) => N317, DATA(25) => N318, DATA(24)
               => N319, DATA(23) => N320, DATA(22) => N321, DATA(21) => N322, 
               DATA(20) => N323, DATA(19) => N324, DATA(18) => N325, DATA(17) 
               => N326, DATA(16) => N327, DATA(15) => N328, DATA(14) => N329, 
               DATA(13) => N330, DATA(12) => N331, DATA(11) => N332, DATA(10) 
               => N333, DATA(9) => N334, DATA(8) => N335, DATA(7) => N336, 
               DATA(6) => N337, DATA(5) => N338, DATA(4) => N339, DATA(3) => 
               N340, DATA(2) => N341, DATA(1) => N342, DATA(0) => N343, 
         -- Connections to port 'DATA2'
         DATA(63) => N507, DATA(62) => N508, DATA(61) => N509, DATA(60) => N510
               , DATA(59) => N511, DATA(58) => N512, DATA(57) => N513, DATA(56)
               => N514, DATA(55) => N515, DATA(54) => N516, DATA(53) => N517, 
               DATA(52) => N518, DATA(51) => N519, DATA(50) => N520, DATA(49) 
               => N521, DATA(48) => N522, DATA(47) => N523, DATA(46) => N524, 
               DATA(45) => N525, DATA(44) => N526, DATA(43) => N527, DATA(42) 
               => N528, DATA(41) => N529, DATA(40) => N530, DATA(39) => N531, 
               DATA(38) => N532, DATA(37) => N533, DATA(36) => N534, DATA(35) 
               => N535, DATA(34) => N536, DATA(33) => N537, DATA(32) => N538, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N13, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N181, 
         -- Connections to port 'Z'
         Z(31) => N604, Z(30) => N603, Z(29) => N602, Z(28) => N601, Z(27) => 
               N600, Z(26) => N599, Z(25) => N598, Z(24) => N597, Z(23) => N596
               , Z(22) => N595, Z(21) => N594, Z(20) => N593, Z(19) => N592, 
               Z(18) => N591, Z(17) => N590, Z(16) => N589, Z(15) => N588, 
               Z(14) => N587, Z(13) => N586, Z(12) => N585, Z(11) => N584, 
               Z(10) => N583, Z(9) => N582, Z(8) => N581, Z(7) => N580, Z(6) =>
               N579, Z(5) => N578, Z(4) => N577, Z(3) => N576, Z(2) => N575, 
               Z(1) => N574, Z(0) => N573 );
   C13938_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic1_port, 
         -- Connections to port 'DATA2'
         DATA(1) => N571, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N13, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N181, 
         -- Connections to port 'Z'
         Z(0) => N605 );
   C13939_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 32 )
      port map(
         -- Connections to port 'DATA1'
         DATA(31) => N474, DATA(30) => N475, DATA(29) => N476, DATA(28) => N477
               , DATA(27) => N478, DATA(26) => N479, DATA(25) => N480, DATA(24)
               => N481, DATA(23) => N482, DATA(22) => N483, DATA(21) => N484, 
               DATA(20) => N485, DATA(19) => N486, DATA(18) => N487, DATA(17) 
               => N488, DATA(16) => N489, DATA(15) => N490, DATA(14) => N491, 
               DATA(13) => N492, DATA(12) => N493, DATA(11) => N494, DATA(10) 
               => N495, DATA(9) => N496, DATA(8) => N497, DATA(7) => N498, 
               DATA(6) => N499, DATA(5) => N500, DATA(4) => N501, DATA(3) => 
               N502, DATA(2) => N503, DATA(1) => N504, DATA(0) => N505, 
         -- Connections to port 'DATA2'
         DATA(63) => N539, DATA(62) => N540, DATA(61) => N541, DATA(60) => N542
               , DATA(59) => N543, DATA(58) => N544, DATA(57) => N545, DATA(56)
               => N546, DATA(55) => N547, DATA(54) => N548, DATA(53) => N549, 
               DATA(52) => N550, DATA(51) => N551, DATA(50) => N552, DATA(49) 
               => N553, DATA(48) => N554, DATA(47) => N555, DATA(46) => N556, 
               DATA(45) => N557, DATA(44) => N558, DATA(43) => N559, DATA(42) 
               => N560, DATA(41) => N561, DATA(40) => N562, DATA(39) => N563, 
               DATA(38) => N564, DATA(37) => N565, DATA(36) => N566, DATA(35) 
               => N567, DATA(34) => N568, DATA(33) => N569, DATA(32) => N570, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N13, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N181, 
         -- Connections to port 'Z'
         Z(31) => N637, Z(30) => N636, Z(29) => N635, Z(28) => N634, Z(27) => 
               N633, Z(26) => N632, Z(25) => N631, Z(24) => N630, Z(23) => N629
               , Z(22) => N628, Z(21) => N627, Z(20) => N626, Z(19) => N625, 
               Z(18) => N624, Z(17) => N623, Z(16) => N622, Z(15) => N621, 
               Z(14) => N620, Z(13) => N619, Z(12) => N618, Z(11) => N617, 
               Z(10) => N616, Z(9) => N615, Z(8) => N614, Z(7) => N613, Z(6) =>
               N612, Z(5) => N611, Z(4) => N610, Z(3) => N609, Z(2) => N608, 
               Z(1) => N607, Z(0) => N606 );
   C13940_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => N572, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N14, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N15, 
         -- Connections to port 'Z'
         Z(0) => N638 );
   B_6 : GTECH_BUF port map( A => ENABLE, Z => N14);
   B_7 : GTECH_BUF port map( A => N179, Z => N15);
   C13941_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => N605, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N14, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N15, 
         -- Connections to port 'Z'
         Z(0) => N639 );
         X_Logic1_port <= '1';
         X_Logic0_port <= '0';
   I_10 : GTECH_NOT port map( A => RESET, Z => N16);
   C13947 : GTECH_AND2 port map( A => ENABLE, B => WR, Z => N17);
   I_11 : GTECH_NOT port map( A => N17, Z => N18);
   I_12 : GTECH_NOT port map( A => ENABLE, Z => N179);
   C14017 : GTECH_AND2 port map( A => RD1_port, B => RD2_port, Z => N180);
   I_13 : GTECH_NOT port map( A => N180, Z => N181);
   I_14 : GTECH_NOT port map( A => ADD_RD1(0), Z => N182);
   I_15 : GTECH_NOT port map( A => ADD_RD1(1), Z => N183);
   C14022 : GTECH_AND2 port map( A => N182, B => N183, Z => N184);
   C14023 : GTECH_AND2 port map( A => N182, B => ADD_RD1(1), Z => N185);
   C14024 : GTECH_AND2 port map( A => ADD_RD1(0), B => N183, Z => N186);
   C14025 : GTECH_AND2 port map( A => ADD_RD1(0), B => ADD_RD1(1), Z => N187);
   I_16 : GTECH_NOT port map( A => ADD_RD1(2), Z => N188);
   C14027 : GTECH_AND2 port map( A => N184, B => N188, Z => N189);
   C14028 : GTECH_AND2 port map( A => N184, B => ADD_RD1(2), Z => N190);
   C14029 : GTECH_AND2 port map( A => N186, B => N188, Z => N191);
   C14030 : GTECH_AND2 port map( A => N186, B => ADD_RD1(2), Z => N192);
   C14031 : GTECH_AND2 port map( A => N185, B => N188, Z => N193);
   C14032 : GTECH_AND2 port map( A => N185, B => ADD_RD1(2), Z => N194);
   C14033 : GTECH_AND2 port map( A => N187, B => N188, Z => N195);
   C14034 : GTECH_AND2 port map( A => N187, B => ADD_RD1(2), Z => N196);
   I_17 : GTECH_NOT port map( A => ADD_RD1(3), Z => N197);
   C14036 : GTECH_AND2 port map( A => N189, B => N197, Z => N198);
   C14037 : GTECH_AND2 port map( A => N189, B => ADD_RD1(3), Z => N199);
   C14038 : GTECH_AND2 port map( A => N191, B => N197, Z => N200);
   C14039 : GTECH_AND2 port map( A => N191, B => ADD_RD1(3), Z => N201);
   C14040 : GTECH_AND2 port map( A => N193, B => N197, Z => N202);
   C14041 : GTECH_AND2 port map( A => N193, B => ADD_RD1(3), Z => N203);
   C14042 : GTECH_AND2 port map( A => N195, B => N197, Z => N204);
   C14043 : GTECH_AND2 port map( A => N195, B => ADD_RD1(3), Z => N205);
   C14044 : GTECH_AND2 port map( A => N190, B => N197, Z => N206);
   C14045 : GTECH_AND2 port map( A => N190, B => ADD_RD1(3), Z => N207);
   C14046 : GTECH_AND2 port map( A => N192, B => N197, Z => N208);
   C14047 : GTECH_AND2 port map( A => N192, B => ADD_RD1(3), Z => N209);
   C14048 : GTECH_AND2 port map( A => N194, B => N197, Z => N210);
   C14049 : GTECH_AND2 port map( A => N194, B => ADD_RD1(3), Z => N211);
   C14050 : GTECH_AND2 port map( A => N196, B => N197, Z => N212);
   C14051 : GTECH_AND2 port map( A => N196, B => ADD_RD1(3), Z => N213);
   I_18 : GTECH_NOT port map( A => ADD_RD1(4), Z => N214);
   C14053 : GTECH_AND2 port map( A => N198, B => N214, Z => N215);
   C14054 : GTECH_AND2 port map( A => N198, B => ADD_RD1(4), Z => N216);
   C14055 : GTECH_AND2 port map( A => N200, B => N214, Z => N217);
   C14056 : GTECH_AND2 port map( A => N200, B => ADD_RD1(4), Z => N218);
   C14057 : GTECH_AND2 port map( A => N202, B => N214, Z => N219);
   C14058 : GTECH_AND2 port map( A => N202, B => ADD_RD1(4), Z => N220);
   C14059 : GTECH_AND2 port map( A => N204, B => N214, Z => N221);
   C14060 : GTECH_AND2 port map( A => N204, B => ADD_RD1(4), Z => N222);
   C14061 : GTECH_AND2 port map( A => N206, B => N214, Z => N223);
   C14062 : GTECH_AND2 port map( A => N206, B => ADD_RD1(4), Z => N224);
   C14063 : GTECH_AND2 port map( A => N208, B => N214, Z => N225);
   C14064 : GTECH_AND2 port map( A => N208, B => ADD_RD1(4), Z => N226);
   C14065 : GTECH_AND2 port map( A => N210, B => N214, Z => N227);
   C14066 : GTECH_AND2 port map( A => N210, B => ADD_RD1(4), Z => N228);
   C14067 : GTECH_AND2 port map( A => N212, B => N214, Z => N229);
   C14068 : GTECH_AND2 port map( A => N212, B => ADD_RD1(4), Z => N230);
   C14069 : GTECH_AND2 port map( A => N199, B => N214, Z => N231);
   C14070 : GTECH_AND2 port map( A => N199, B => ADD_RD1(4), Z => N232);
   C14071 : GTECH_AND2 port map( A => N201, B => N214, Z => N233);
   C14072 : GTECH_AND2 port map( A => N201, B => ADD_RD1(4), Z => N234);
   C14073 : GTECH_AND2 port map( A => N203, B => N214, Z => N235);
   C14074 : GTECH_AND2 port map( A => N203, B => ADD_RD1(4), Z => N236);
   C14075 : GTECH_AND2 port map( A => N205, B => N214, Z => N237);
   C14076 : GTECH_AND2 port map( A => N205, B => ADD_RD1(4), Z => N238);
   C14077 : GTECH_AND2 port map( A => N207, B => N214, Z => N239);
   C14078 : GTECH_AND2 port map( A => N207, B => ADD_RD1(4), Z => N240);
   C14079 : GTECH_AND2 port map( A => N209, B => N214, Z => N241);
   C14080 : GTECH_AND2 port map( A => N209, B => ADD_RD1(4), Z => N242);
   C14081 : GTECH_AND2 port map( A => N211, B => N214, Z => N243);
   C14082 : GTECH_AND2 port map( A => N211, B => ADD_RD1(4), Z => N244);
   C14083 : GTECH_AND2 port map( A => N213, B => N214, Z => N245);
   C14084 : GTECH_AND2 port map( A => N213, B => ADD_RD1(4), Z => N246);
   I_19 : GTECH_NOT port map( A => ADD_RD1(5), Z => N247);
   C14086 : GTECH_AND2 port map( A => N215, B => N247, Z => N248);
   C14087 : GTECH_AND2 port map( A => N215, B => ADD_RD1(5), Z => N249);
   C14088 : GTECH_AND2 port map( A => N217, B => N247, Z => N250);
   C14089 : GTECH_AND2 port map( A => N217, B => ADD_RD1(5), Z => N251);
   C14090 : GTECH_AND2 port map( A => N219, B => N247, Z => N252);
   C14091 : GTECH_AND2 port map( A => N219, B => ADD_RD1(5), Z => N253);
   C14092 : GTECH_AND2 port map( A => N221, B => N247, Z => N254);
   C14093 : GTECH_AND2 port map( A => N221, B => ADD_RD1(5), Z => N255);
   C14094 : GTECH_AND2 port map( A => N223, B => N247, Z => N256);
   C14095 : GTECH_AND2 port map( A => N223, B => ADD_RD1(5), Z => N257);
   C14096 : GTECH_AND2 port map( A => N225, B => N247, Z => N258);
   C14097 : GTECH_AND2 port map( A => N225, B => ADD_RD1(5), Z => N259);
   C14098 : GTECH_AND2 port map( A => N227, B => N247, Z => N260);
   C14099 : GTECH_AND2 port map( A => N227, B => ADD_RD1(5), Z => N261);
   C14100 : GTECH_AND2 port map( A => N229, B => N247, Z => N262);
   C14101 : GTECH_AND2 port map( A => N229, B => ADD_RD1(5), Z => N263);
   C14102 : GTECH_AND2 port map( A => N231, B => N247, Z => N264);
   C14103 : GTECH_AND2 port map( A => N231, B => ADD_RD1(5), Z => N265);
   C14104 : GTECH_AND2 port map( A => N233, B => N247, Z => N266);
   C14105 : GTECH_AND2 port map( A => N233, B => ADD_RD1(5), Z => N267);
   C14106 : GTECH_AND2 port map( A => N235, B => N247, Z => N268);
   C14107 : GTECH_AND2 port map( A => N235, B => ADD_RD1(5), Z => N269);
   C14108 : GTECH_AND2 port map( A => N237, B => N247, Z => N270);
   C14109 : GTECH_AND2 port map( A => N237, B => ADD_RD1(5), Z => N271);
   C14110 : GTECH_AND2 port map( A => N239, B => N247, Z => N272);
   C14111 : GTECH_AND2 port map( A => N239, B => ADD_RD1(5), Z => N273);
   C14112 : GTECH_AND2 port map( A => N241, B => N247, Z => N274);
   C14113 : GTECH_AND2 port map( A => N241, B => ADD_RD1(5), Z => N275);
   C14114 : GTECH_AND2 port map( A => N243, B => N247, Z => N276);
   C14115 : GTECH_AND2 port map( A => N243, B => ADD_RD1(5), Z => N277);
   C14116 : GTECH_AND2 port map( A => N245, B => N247, Z => N278);
   C14117 : GTECH_AND2 port map( A => N245, B => ADD_RD1(5), Z => N279);
   C14118 : GTECH_AND2 port map( A => N216, B => N247, Z => N280);
   C14119 : GTECH_AND2 port map( A => N216, B => ADD_RD1(5), Z => N281);
   C14120 : GTECH_AND2 port map( A => N218, B => N247, Z => N282);
   C14121 : GTECH_AND2 port map( A => N218, B => ADD_RD1(5), Z => N283);
   C14122 : GTECH_AND2 port map( A => N220, B => N247, Z => N284);
   C14123 : GTECH_AND2 port map( A => N220, B => ADD_RD1(5), Z => N285);
   C14124 : GTECH_AND2 port map( A => N222, B => N247, Z => N286);
   C14125 : GTECH_AND2 port map( A => N222, B => ADD_RD1(5), Z => N287);
   C14126 : GTECH_AND2 port map( A => N224, B => N247, Z => N288);
   C14127 : GTECH_AND2 port map( A => N224, B => ADD_RD1(5), Z => N289);
   C14128 : GTECH_AND2 port map( A => N226, B => N247, Z => N290);
   C14129 : GTECH_AND2 port map( A => N226, B => ADD_RD1(5), Z => N291);
   C14130 : GTECH_AND2 port map( A => N228, B => N247, Z => N292);
   C14131 : GTECH_AND2 port map( A => N228, B => ADD_RD1(5), Z => N293);
   C14132 : GTECH_AND2 port map( A => N230, B => N247, Z => N294);
   C14133 : GTECH_AND2 port map( A => N230, B => ADD_RD1(5), Z => N295);
   C14134 : GTECH_AND2 port map( A => N232, B => N247, Z => N296);
   C14135 : GTECH_AND2 port map( A => N232, B => ADD_RD1(5), Z => N297);
   C14136 : GTECH_AND2 port map( A => N234, B => N247, Z => N298);
   C14137 : GTECH_AND2 port map( A => N234, B => ADD_RD1(5), Z => N299);
   C14138 : GTECH_AND2 port map( A => N236, B => N247, Z => N300);
   C14139 : GTECH_AND2 port map( A => N236, B => ADD_RD1(5), Z => N301);
   C14140 : GTECH_AND2 port map( A => N238, B => N247, Z => N302);
   C14141 : GTECH_AND2 port map( A => N238, B => ADD_RD1(5), Z => N303);
   C14142 : GTECH_AND2 port map( A => N240, B => N247, Z => N304);
   C14143 : GTECH_AND2 port map( A => N240, B => ADD_RD1(5), Z => N305);
   C14144 : GTECH_AND2 port map( A => N242, B => N247, Z => N306);
   C14145 : GTECH_AND2 port map( A => N242, B => ADD_RD1(5), Z => N307);
   C14146 : GTECH_AND2 port map( A => N244, B => N247, Z => N308);
   C14147 : GTECH_AND2 port map( A => N244, B => ADD_RD1(5), Z => N309);
   C14148 : GTECH_AND2 port map( A => N246, B => N247, Z => N310);
   C14149 : GTECH_AND2 port map( A => N246, B => ADD_RD1(5), Z => N311);
   I_20 : GTECH_NOT port map( A => ADD_RD2(0), Z => N344);
   I_21 : GTECH_NOT port map( A => ADD_RD2(1), Z => N345);
   C14152 : GTECH_AND2 port map( A => N344, B => N345, Z => N346);
   C14153 : GTECH_AND2 port map( A => N344, B => ADD_RD2(1), Z => N347);
   C14154 : GTECH_AND2 port map( A => ADD_RD2(0), B => N345, Z => N348);
   C14155 : GTECH_AND2 port map( A => ADD_RD2(0), B => ADD_RD2(1), Z => N349);
   I_22 : GTECH_NOT port map( A => ADD_RD2(2), Z => N350);
   C14157 : GTECH_AND2 port map( A => N346, B => N350, Z => N351);
   C14158 : GTECH_AND2 port map( A => N346, B => ADD_RD2(2), Z => N352);
   C14159 : GTECH_AND2 port map( A => N348, B => N350, Z => N353);
   C14160 : GTECH_AND2 port map( A => N348, B => ADD_RD2(2), Z => N354);
   C14161 : GTECH_AND2 port map( A => N347, B => N350, Z => N355);
   C14162 : GTECH_AND2 port map( A => N347, B => ADD_RD2(2), Z => N356);
   C14163 : GTECH_AND2 port map( A => N349, B => N350, Z => N357);
   C14164 : GTECH_AND2 port map( A => N349, B => ADD_RD2(2), Z => N358);
   I_23 : GTECH_NOT port map( A => ADD_RD2(3), Z => N359);
   C14166 : GTECH_AND2 port map( A => N351, B => N359, Z => N360);
   C14167 : GTECH_AND2 port map( A => N351, B => ADD_RD2(3), Z => N361);
   C14168 : GTECH_AND2 port map( A => N353, B => N359, Z => N362);
   C14169 : GTECH_AND2 port map( A => N353, B => ADD_RD2(3), Z => N363);
   C14170 : GTECH_AND2 port map( A => N355, B => N359, Z => N364);
   C14171 : GTECH_AND2 port map( A => N355, B => ADD_RD2(3), Z => N365);
   C14172 : GTECH_AND2 port map( A => N357, B => N359, Z => N366);
   C14173 : GTECH_AND2 port map( A => N357, B => ADD_RD2(3), Z => N367);
   C14174 : GTECH_AND2 port map( A => N352, B => N359, Z => N368);
   C14175 : GTECH_AND2 port map( A => N352, B => ADD_RD2(3), Z => N369);
   C14176 : GTECH_AND2 port map( A => N354, B => N359, Z => N370);
   C14177 : GTECH_AND2 port map( A => N354, B => ADD_RD2(3), Z => N371);
   C14178 : GTECH_AND2 port map( A => N356, B => N359, Z => N372);
   C14179 : GTECH_AND2 port map( A => N356, B => ADD_RD2(3), Z => N373);
   C14180 : GTECH_AND2 port map( A => N358, B => N359, Z => N374);
   C14181 : GTECH_AND2 port map( A => N358, B => ADD_RD2(3), Z => N375);
   I_24 : GTECH_NOT port map( A => ADD_RD2(4), Z => N376);
   C14183 : GTECH_AND2 port map( A => N360, B => N376, Z => N377);
   C14184 : GTECH_AND2 port map( A => N360, B => ADD_RD2(4), Z => N378);
   C14185 : GTECH_AND2 port map( A => N362, B => N376, Z => N379);
   C14186 : GTECH_AND2 port map( A => N362, B => ADD_RD2(4), Z => N380);
   C14187 : GTECH_AND2 port map( A => N364, B => N376, Z => N381);
   C14188 : GTECH_AND2 port map( A => N364, B => ADD_RD2(4), Z => N382);
   C14189 : GTECH_AND2 port map( A => N366, B => N376, Z => N383);
   C14190 : GTECH_AND2 port map( A => N366, B => ADD_RD2(4), Z => N384);
   C14191 : GTECH_AND2 port map( A => N368, B => N376, Z => N385);
   C14192 : GTECH_AND2 port map( A => N368, B => ADD_RD2(4), Z => N386);
   C14193 : GTECH_AND2 port map( A => N370, B => N376, Z => N387);
   C14194 : GTECH_AND2 port map( A => N370, B => ADD_RD2(4), Z => N388);
   C14195 : GTECH_AND2 port map( A => N372, B => N376, Z => N389);
   C14196 : GTECH_AND2 port map( A => N372, B => ADD_RD2(4), Z => N390);
   C14197 : GTECH_AND2 port map( A => N374, B => N376, Z => N391);
   C14198 : GTECH_AND2 port map( A => N374, B => ADD_RD2(4), Z => N392);
   C14199 : GTECH_AND2 port map( A => N361, B => N376, Z => N393);
   C14200 : GTECH_AND2 port map( A => N361, B => ADD_RD2(4), Z => N394);
   C14201 : GTECH_AND2 port map( A => N363, B => N376, Z => N395);
   C14202 : GTECH_AND2 port map( A => N363, B => ADD_RD2(4), Z => N396);
   C14203 : GTECH_AND2 port map( A => N365, B => N376, Z => N397);
   C14204 : GTECH_AND2 port map( A => N365, B => ADD_RD2(4), Z => N398);
   C14205 : GTECH_AND2 port map( A => N367, B => N376, Z => N399);
   C14206 : GTECH_AND2 port map( A => N367, B => ADD_RD2(4), Z => N400);
   C14207 : GTECH_AND2 port map( A => N369, B => N376, Z => N401);
   C14208 : GTECH_AND2 port map( A => N369, B => ADD_RD2(4), Z => N402);
   C14209 : GTECH_AND2 port map( A => N371, B => N376, Z => N403);
   C14210 : GTECH_AND2 port map( A => N371, B => ADD_RD2(4), Z => N404);
   C14211 : GTECH_AND2 port map( A => N373, B => N376, Z => N405);
   C14212 : GTECH_AND2 port map( A => N373, B => ADD_RD2(4), Z => N406);
   C14213 : GTECH_AND2 port map( A => N375, B => N376, Z => N407);
   C14214 : GTECH_AND2 port map( A => N375, B => ADD_RD2(4), Z => N408);
   I_25 : GTECH_NOT port map( A => ADD_RD2(5), Z => N409);
   C14216 : GTECH_AND2 port map( A => N377, B => N409, Z => N410);
   C14217 : GTECH_AND2 port map( A => N377, B => ADD_RD2(5), Z => N411);
   C14218 : GTECH_AND2 port map( A => N379, B => N409, Z => N412);
   C14219 : GTECH_AND2 port map( A => N379, B => ADD_RD2(5), Z => N413);
   C14220 : GTECH_AND2 port map( A => N381, B => N409, Z => N414);
   C14221 : GTECH_AND2 port map( A => N381, B => ADD_RD2(5), Z => N415);
   C14222 : GTECH_AND2 port map( A => N383, B => N409, Z => N416);
   C14223 : GTECH_AND2 port map( A => N383, B => ADD_RD2(5), Z => N417);
   C14224 : GTECH_AND2 port map( A => N385, B => N409, Z => N418);
   C14225 : GTECH_AND2 port map( A => N385, B => ADD_RD2(5), Z => N419);
   C14226 : GTECH_AND2 port map( A => N387, B => N409, Z => N420);
   C14227 : GTECH_AND2 port map( A => N387, B => ADD_RD2(5), Z => N421);
   C14228 : GTECH_AND2 port map( A => N389, B => N409, Z => N422);
   C14229 : GTECH_AND2 port map( A => N389, B => ADD_RD2(5), Z => N423);
   C14230 : GTECH_AND2 port map( A => N391, B => N409, Z => N424);
   C14231 : GTECH_AND2 port map( A => N391, B => ADD_RD2(5), Z => N425);
   C14232 : GTECH_AND2 port map( A => N393, B => N409, Z => N426);
   C14233 : GTECH_AND2 port map( A => N393, B => ADD_RD2(5), Z => N427);
   C14234 : GTECH_AND2 port map( A => N395, B => N409, Z => N428);
   C14235 : GTECH_AND2 port map( A => N395, B => ADD_RD2(5), Z => N429);
   C14236 : GTECH_AND2 port map( A => N397, B => N409, Z => N430);
   C14237 : GTECH_AND2 port map( A => N397, B => ADD_RD2(5), Z => N431);
   C14238 : GTECH_AND2 port map( A => N399, B => N409, Z => N432);
   C14239 : GTECH_AND2 port map( A => N399, B => ADD_RD2(5), Z => N433);
   C14240 : GTECH_AND2 port map( A => N401, B => N409, Z => N434);
   C14241 : GTECH_AND2 port map( A => N401, B => ADD_RD2(5), Z => N435);
   C14242 : GTECH_AND2 port map( A => N403, B => N409, Z => N436);
   C14243 : GTECH_AND2 port map( A => N403, B => ADD_RD2(5), Z => N437);
   C14244 : GTECH_AND2 port map( A => N405, B => N409, Z => N438);
   C14245 : GTECH_AND2 port map( A => N405, B => ADD_RD2(5), Z => N439);
   C14246 : GTECH_AND2 port map( A => N407, B => N409, Z => N440);
   C14247 : GTECH_AND2 port map( A => N407, B => ADD_RD2(5), Z => N441);
   C14248 : GTECH_AND2 port map( A => N378, B => N409, Z => N442);
   C14249 : GTECH_AND2 port map( A => N378, B => ADD_RD2(5), Z => N443);
   C14250 : GTECH_AND2 port map( A => N380, B => N409, Z => N444);
   C14251 : GTECH_AND2 port map( A => N380, B => ADD_RD2(5), Z => N445);
   C14252 : GTECH_AND2 port map( A => N382, B => N409, Z => N446);
   C14253 : GTECH_AND2 port map( A => N382, B => ADD_RD2(5), Z => N447);
   C14254 : GTECH_AND2 port map( A => N384, B => N409, Z => N448);
   C14255 : GTECH_AND2 port map( A => N384, B => ADD_RD2(5), Z => N449);
   C14256 : GTECH_AND2 port map( A => N386, B => N409, Z => N450);
   C14257 : GTECH_AND2 port map( A => N386, B => ADD_RD2(5), Z => N451);
   C14258 : GTECH_AND2 port map( A => N388, B => N409, Z => N452);
   C14259 : GTECH_AND2 port map( A => N388, B => ADD_RD2(5), Z => N453);
   C14260 : GTECH_AND2 port map( A => N390, B => N409, Z => N454);
   C14261 : GTECH_AND2 port map( A => N390, B => ADD_RD2(5), Z => N455);
   C14262 : GTECH_AND2 port map( A => N392, B => N409, Z => N456);
   C14263 : GTECH_AND2 port map( A => N392, B => ADD_RD2(5), Z => N457);
   C14264 : GTECH_AND2 port map( A => N394, B => N409, Z => N458);
   C14265 : GTECH_AND2 port map( A => N394, B => ADD_RD2(5), Z => N459);
   C14266 : GTECH_AND2 port map( A => N396, B => N409, Z => N460);
   C14267 : GTECH_AND2 port map( A => N396, B => ADD_RD2(5), Z => N461);
   C14268 : GTECH_AND2 port map( A => N398, B => N409, Z => N462);
   C14269 : GTECH_AND2 port map( A => N398, B => ADD_RD2(5), Z => N463);
   C14270 : GTECH_AND2 port map( A => N400, B => N409, Z => N464);
   C14271 : GTECH_AND2 port map( A => N400, B => ADD_RD2(5), Z => N465);
   C14272 : GTECH_AND2 port map( A => N402, B => N409, Z => N466);
   C14273 : GTECH_AND2 port map( A => N402, B => ADD_RD2(5), Z => N467);
   C14274 : GTECH_AND2 port map( A => N404, B => N409, Z => N468);
   C14275 : GTECH_AND2 port map( A => N404, B => ADD_RD2(5), Z => N469);
   C14276 : GTECH_AND2 port map( A => N406, B => N409, Z => N470);
   C14277 : GTECH_AND2 port map( A => N406, B => ADD_RD2(5), Z => N471);
   C14278 : GTECH_AND2 port map( A => N408, B => N409, Z => N472);
   C14279 : GTECH_AND2 port map( A => N408, B => ADD_RD2(5), Z => N473);
   I_26 : GTECH_NOT port map( A => RD1_port, Z => N506);

end SYN_Beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_topLevel_1.all;

entity RMU_M8_N8_F3_VIRTUAL_ADDR_SIZE5_PHY_ADDR_SIZE6 is

   port( CALL, RET : in std_logic;  STALL : out std_logic;  READ1, READ2, WRITE
         : in std_logic;  RD1, RD2, WR : out std_logic;  ENABLE, RST, CLK : in 
         std_logic;  SPILL, FILL : out std_logic;  ACK : in std_logic;  
         PHY_ADDRESS1, PHY_ADDRESS2, PHY_ADDRESS3 : out std_logic_vector (5 
         downto 0);  VIRTUAL_ADDRESS1, VIRTUAL_ADDRESS2, VIRTUAL_ADDRESS3 : in 
         std_logic_vector (4 downto 0));

end RMU_M8_N8_F3_VIRTUAL_ADDR_SIZE5_PHY_ADDR_SIZE6;

architecture SYN_HLSM of RMU_M8_N8_F3_VIRTUAL_ADDR_SIZE5_PHY_ADDR_SIZE6 is

   component GTECH_AND2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component GTECH_NOT
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component GTECH_BUF
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component GTECH_OR2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component GTECH_OR4
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component GTECH_OR3
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
      generic ( ac_as_q, ac_as_qn, sc_ss_q : integer );
      port(
         clear, preset, enable, data_in, synch_clear, synch_preset, 
            synch_toggle, synch_enable, next_state, clocked_on : in std_logic;
         Q, QN : buffer std_logic
      );
   end component;
   
   component MOD_UNS_OP
      generic( A_width, B_width, REMAINDER_width : integer );
      port( A : in std_logic_vector(A_width - 1 downto 0); B : in 
            std_logic_vector(B_width - 1 downto 0); REMAINDER : out 
            std_logic_vector(REMAINDER_width - 1 downto 0) );
   end component;
   
   signal N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
      N16, N17, N18, X_Logic1_port, X_Logic0_port, CALL_port, RET_port, 
      STALL_port, READ1_port, READ2_port, WRITE_port, RD1_port, RD2_port, 
      WR_port, ENABLE_port, CLK_port, SPILL_port, FILL_port, 
      PHY_ADDRESS1_5_port, PHY_ADDRESS1_4_port, PHY_ADDRESS1_3_port, 
      PHY_ADDRESS1_2_port, PHY_ADDRESS1_1_port, PHY_ADDRESS1_0_port, 
      PHY_ADDRESS2_5_port, PHY_ADDRESS2_4_port, PHY_ADDRESS2_3_port, 
      PHY_ADDRESS2_2_port, PHY_ADDRESS2_1_port, PHY_ADDRESS2_0_port, 
      PHY_ADDRESS3_5_port, PHY_ADDRESS3_4_port, PHY_ADDRESS3_3_port, 
      PHY_ADDRESS3_2_port, PHY_ADDRESS3_1_port, PHY_ADDRESS3_0_port, 
      VIRTUAL_ADDRESS1_4_port, VIRTUAL_ADDRESS1_3_port, VIRTUAL_ADDRESS1_2_port
      , VIRTUAL_ADDRESS1_1_port, VIRTUAL_ADDRESS1_0_port, 
      VIRTUAL_ADDRESS2_4_port, VIRTUAL_ADDRESS2_3_port, VIRTUAL_ADDRESS2_2_port
      , VIRTUAL_ADDRESS2_1_port, VIRTUAL_ADDRESS2_0_port, 
      VIRTUAL_ADDRESS3_4_port, VIRTUAL_ADDRESS3_3_port, VIRTUAL_ADDRESS3_2_port
      , VIRTUAL_ADDRESS3_1_port, VIRTUAL_ADDRESS3_0_port, N19, 
      curr_state_2_port, curr_state_1_port, curr_state_0_port, 
      curr_CANSAVE_1_port, curr_CANSAVE_0_port, next_state_2_port, 
      next_state_1_port, next_state_0_port, next_CWP_6_port, next_CWP_5_port, 
      next_CWP_4_port, next_CWP_3_port, next_CWP_2_port, next_CWP_1_port, 
      next_CWP_0_port, next_SWP_6_port, next_SWP_5_port, next_SWP_4_port, 
      next_SWP_3_port, next_SWP_2_port, next_SWP_1_port, next_SWP_0_port, 
      next_RESTORE_6_port, next_RESTORE_5_port, next_RESTORE_4_port, 
      next_RESTORE_3_port, next_RESTORE_2_port, next_RESTORE_1_port, 
      next_RESTORE_0_port, next_CANSAVE_1_port, next_CANSAVE_0_port, N20, N21, 
      N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36
      , N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, net30, N48, 
      net31, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, 
      N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73, net33, N74, 
      net34, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, 
      N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, net36, N100, 
      net37, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110, N111, 
      N112, N113, N114, N115, N116, N117, N118, N119, N120, N121, N122, N123, 
      N124, N125, N126, N127, N128, N129, N130, N131, N132, N133, N134, N135, 
      N136, N137, N138, N139, N140, N141, N142, N143, N144, N145, N146, N147, 
      N148, N149, N150, N151, N152, N153, N154, N155, N156, N157, N158, N159, 
      N160, N161, N162, N163, N164, N165, N166, N167, N168, N169, N170, N171, 
      N172, N173, N174, N175, N176, N177, N178, N179, N180, N181, N182, N183, 
      N184, N185, N186, N187, N188, N189, N190, N191, N192, N193, N194, N195, 
      N196, N197, N198, N199, N200, N201, N202, N203, N204, N205, N206, N207, 
      N208, N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, 
      N220, N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231, 
      N232, N233, N234, N235, N236, N237, N238, N239, N240, N241, N242, N243, 
      N244, N245, N246, N247, N248, N249, N250, N251, N252, N253, N254, N255, 
      N256, N257, N258, N259, N260, N261, N262, N263, N264, N265, N266, N267, 
      N268, N269, N270, N271, N272, N273, N274, N275, N276, N277, N278, N279, 
      N280, N281, N282, N283, N284, N285, N286, N287, N288, N289, n_3112, 
      n_3113, n_3114, n_3115, n_3116, n_3117, n_3118, n_3119, n_3120, n_3121, 
      n_3122, n_3123, n_3124, n_3125, n_3126, n_3127, n_3128, n_3129, n_3130, 
      n_3131, n_3132, n_3133, n_3134, n_3135, n_3136, n_3137, n_3138, n_3139, 
      n_3140, n_3141, n_3142, n_3143, n_3144, n_3145, n_3146, n_3147, n_3148, 
      n_3149, n_3150, n_3151, n_3152, n_3153, n_3154, n_3155, n_3156, n_3157, 
      n_3158, n_3159, n_3160, n_3161, n_3162, n_3163, n_3164, n_3165, n_3166, 
      n_3167, n_3168, n_3169, n_3170, n_3171, n_3172, n_3173, n_3174, n_3175, 
      n_3176, n_3177, n_3178, n_3179, n_3180, n_3181, n_3182, n_3183, n_3184, 
      n_3185, n_3186, n_3187, n_3188, n_3189, n_3190, n_3191, n_3192, n_3193, 
      n_3194, n_3195, n_3196, n_3197, n_3198, n_3199, n_3200, n_3201, n_3202, 
      n_3203, n_3204, n_3205, n_3206, n_3207, n_3208, n_3209, n_3210, n_3211, 
      n_3212, n_3213, n_3214, n_3215, n_3216, n_3217, n_3218, n_3219, n_3220, 
      n_3221, n_3222, n_3223, n_3224, n_3225, n_3226, n_3227, n_3228, n_3229, 
      n_3230, n_3231, n_3232, n_3233, n_3234, n_3235, n_3236, n_3237, n_3238, 
      n_3239, n_3240, n_3241, n_3242, n_3243, n_3244, n_3245, n_3246, n_3247, 
      n_3248, n_3249, n_3250, n_3251, n_3252, n_3253, n_3254, n_3255, n_3256, 
      n_3257, n_3258, n_3259, n_3260, n_3261, n_3262, n_3263, n_3264, n_3265, 
      n_3266, n_3267, n_3268, n_3269, n_3270, n_3271, n_3272, n_3273, n_3274, 
      n_3275, n_3276, n_3277, n_3278, n_3279, n_3280, n_3281, n_3282, n_3283, 
      n_3284, n_3285, n_3286, n_3287, n_3288, n_3289, n_3290, n_3291, n_3292, 
      n_3293, n_3294, n_3295, n_3296, n_3297, n_3298, n_3299, n_3300, n_3301, 
      n_3302, n_3303, n_3304, n_3305, n_3306, n_3307, n_3308, n_3309, n_3310, 
      n_3311, n_3312, n_3313, n_3314, n_3315, n_3316, n_3317, n_3318, n_3319, 
      n_3320, n_3321, n_3322, n_3323, n_3324, n_3325, n_3326, n_3327, n_3328, 
      n_3329, n_3330, n_3331, n_3332, n_3333, n_3334, n_3335, n_3336, n_3337, 
      n_3338, n_3339, n_3340, n_3341, n_3342, n_3343, n_3344, n_3345, n_3346, 
      n_3347, n_3348, n_3349, n_3350, n_3351, n_3352, n_3353, n_3354, n_3355, 
      n_3356, n_3357, n_3358, n_3359, n_3360, n_3361, n_3362 : std_logic;

begin
   CALL_port <= CALL;
   RET_port <= RET;
   STALL <= STALL_port;
   READ1_port <= READ1;
   READ2_port <= READ2;
   WRITE_port <= WRITE;
   RD1 <= RD1_port;
   RD2 <= RD2_port;
   WR <= WR_port;
   ENABLE_port <= ENABLE;
   CLK_port <= CLK;
   SPILL <= SPILL_port;
   FILL <= FILL_port;
   PHY_ADDRESS1 <= ( PHY_ADDRESS1_5_port, PHY_ADDRESS1_4_port, 
      PHY_ADDRESS1_3_port, PHY_ADDRESS1_2_port, PHY_ADDRESS1_1_port, 
      PHY_ADDRESS1_0_port );
   PHY_ADDRESS2 <= ( PHY_ADDRESS2_5_port, PHY_ADDRESS2_4_port, 
      PHY_ADDRESS2_3_port, PHY_ADDRESS2_2_port, PHY_ADDRESS2_1_port, 
      PHY_ADDRESS2_0_port );
   PHY_ADDRESS3 <= ( PHY_ADDRESS3_5_port, PHY_ADDRESS3_4_port, 
      PHY_ADDRESS3_3_port, PHY_ADDRESS3_2_port, PHY_ADDRESS3_1_port, 
      PHY_ADDRESS3_0_port );
   ( VIRTUAL_ADDRESS1_4_port, VIRTUAL_ADDRESS1_3_port, VIRTUAL_ADDRESS1_2_port,
      VIRTUAL_ADDRESS1_1_port, VIRTUAL_ADDRESS1_0_port ) <= VIRTUAL_ADDRESS1;
   ( VIRTUAL_ADDRESS2_4_port, VIRTUAL_ADDRESS2_3_port, VIRTUAL_ADDRESS2_2_port,
      VIRTUAL_ADDRESS2_1_port, VIRTUAL_ADDRESS2_0_port ) <= VIRTUAL_ADDRESS2;
   ( VIRTUAL_ADDRESS3_4_port, VIRTUAL_ADDRESS3_3_port, VIRTUAL_ADDRESS3_2_port,
      VIRTUAL_ADDRESS3_1_port, VIRTUAL_ADDRESS3_0_port ) <= VIRTUAL_ADDRESS3;
   
   curr_CANSAVE_reg_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N20, next_state => N46, 
               clocked_on => CLK_port, Q => curr_CANSAVE_1_port, QN => n_3112);
   curr_CANSAVE_reg_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N20, next_state => N45, 
               clocked_on => CLK_port, Q => curr_CANSAVE_0_port, QN => n_3113);
   curr_state_reg_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N20, next_state => N23, 
               clocked_on => CLK_port, Q => curr_state_2_port, QN => n_3114);
   curr_state_reg_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N20, next_state => N22, 
               clocked_on => CLK_port, Q => curr_state_1_port, QN => n_3115);
   curr_state_reg_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N20, next_state => N21, 
               clocked_on => CLK_port, Q => curr_state_0_port, QN => n_3116);
   curr_CWP_reg_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N20, next_state => N30, 
               clocked_on => CLK_port, Q => N272, QN => n_3117);
   curr_CWP_reg_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N20, next_state => N29, 
               clocked_on => CLK_port, Q => N273, QN => n_3118);
   curr_CWP_reg_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N20, next_state => N28, 
               clocked_on => CLK_port, Q => N274, QN => n_3119);
   curr_CWP_reg_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N20, next_state => N27, 
               clocked_on => CLK_port, Q => N275, QN => n_3120);
   curr_CWP_reg_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N20, next_state => N26, 
               clocked_on => CLK_port, Q => N276, QN => n_3121);
   curr_CWP_reg_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N20, next_state => N25, 
               clocked_on => CLK_port, Q => N277, QN => n_3122);
   curr_CWP_reg_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N20, next_state => N24, 
               clocked_on => CLK_port, Q => N278, QN => n_3123);
   curr_SWP_reg_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N20, next_state => N37, 
               clocked_on => CLK_port, Q => N280, QN => n_3124);
   curr_SWP_reg_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N20, next_state => N36, 
               clocked_on => CLK_port, Q => N281, QN => n_3125);
   curr_SWP_reg_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N20, next_state => N35, 
               clocked_on => CLK_port, Q => N282, QN => n_3126);
   curr_SWP_reg_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N20, next_state => N34, 
               clocked_on => CLK_port, Q => N283, QN => n_3127);
   curr_SWP_reg_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N20, next_state => N33, 
               clocked_on => CLK_port, Q => N284, QN => n_3128);
   curr_SWP_reg_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N20, next_state => N32, 
               clocked_on => CLK_port, Q => N285, QN => n_3129);
   curr_SWP_reg_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N20, next_state => N31, 
               clocked_on => CLK_port, Q => N286, QN => n_3130);
   curr_RESTORE_reg_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N20, next_state => N44, 
               clocked_on => CLK_port, Q => N265, QN => n_3131);
   curr_RESTORE_reg_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N20, next_state => N43, 
               clocked_on => CLK_port, Q => N266, QN => n_3132);
   curr_RESTORE_reg_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N20, next_state => N42, 
               clocked_on => CLK_port, Q => N267, QN => n_3133);
   curr_RESTORE_reg_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N20, next_state => N41, 
               clocked_on => CLK_port, Q => N268, QN => n_3134);
   curr_RESTORE_reg_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N20, next_state => N40, 
               clocked_on => CLK_port, Q => N269, QN => n_3135);
   curr_RESTORE_reg_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N20, next_state => N39, 
               clocked_on => CLK_port, Q => N270, QN => n_3136);
   curr_RESTORE_reg_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N20, next_state => N38, 
               clocked_on => CLK_port, Q => N271, QN => n_3137);
   lt_85 : process ( X_Logic0_port, VIRTUAL_ADDRESS1_4_port, 
         VIRTUAL_ADDRESS1_3_port, VIRTUAL_ADDRESS1_2_port, 
         VIRTUAL_ADDRESS1_1_port, VIRTUAL_ADDRESS1_0_port, X_Logic1_port )
      variable A : SIGNED( 5 downto 0 );
      variable B : SIGNED( 4 downto 0 );
      variable Z : SIGNED( 0 downto 0 );
   begin
      A := ( X_Logic0_port, VIRTUAL_ADDRESS1_4_port, VIRTUAL_ADDRESS1_3_port, 
            VIRTUAL_ADDRESS1_2_port, VIRTUAL_ADDRESS1_1_port, 
            VIRTUAL_ADDRESS1_0_port );
      B := ( X_Logic0_port, X_Logic1_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port );
      if ( A < B ) then
         Z := ( others => '1' );
      else
         Z := ( others => '0' );
      end if;
      ( 0 => N47 ) <= Z;
   end process;
   
   mod_91 : MOD_UNS_OP
      generic map ( A_width => 6, B_width => 31, REMAINDER_width => 31 )
      port map(
         -- Connections to port 'A'
         A(5) => N66, A(4) => N65, A(3) => N64, A(2) => N63, A(1) => N62, A(0) 
               => N61, 
         -- Connections to port 'B'
         B(30) => X_Logic0_port, B(29) => X_Logic0_port, B(28) => X_Logic0_port
               , B(27) => X_Logic0_port, B(26) => X_Logic0_port, B(25) => 
               X_Logic0_port, B(24) => X_Logic0_port, B(23) => X_Logic0_port, 
               B(22) => X_Logic0_port, B(21) => X_Logic0_port, B(20) => 
               X_Logic0_port, B(19) => X_Logic0_port, B(18) => X_Logic0_port, 
               B(17) => X_Logic0_port, B(16) => X_Logic0_port, B(15) => 
               X_Logic0_port, B(14) => X_Logic0_port, B(13) => X_Logic0_port, 
               B(12) => X_Logic0_port, B(11) => X_Logic0_port, B(10) => 
               X_Logic0_port, B(9) => X_Logic0_port, B(8) => X_Logic0_port, 
               B(7) => X_Logic0_port, B(6) => X_Logic0_port, B(5) => 
               X_Logic1_port, B(4) => X_Logic1_port, B(3) => X_Logic1_port, 
               B(2) => X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
               X_Logic0_port, 
         -- Connections to port 'REMAINDER'
         REMAINDER(30) => n_3138, REMAINDER(29) => n_3139, REMAINDER(28) => 
               n_3140, REMAINDER(27) => n_3141, REMAINDER(26) => n_3142, 
               REMAINDER(25) => n_3143, REMAINDER(24) => n_3144, REMAINDER(23) 
               => n_3145, REMAINDER(22) => n_3146, REMAINDER(21) => n_3147, 
               REMAINDER(20) => n_3148, REMAINDER(19) => n_3149, REMAINDER(18) 
               => n_3150, REMAINDER(17) => n_3151, REMAINDER(16) => n_3152, 
               REMAINDER(15) => n_3153, REMAINDER(14) => n_3154, REMAINDER(13) 
               => n_3155, REMAINDER(12) => n_3156, REMAINDER(11) => n_3157, 
               REMAINDER(10) => n_3158, REMAINDER(9) => n_3159, REMAINDER(8) =>
               n_3160, REMAINDER(7) => n_3161, REMAINDER(6) => n_3162, 
               REMAINDER(5) => N72, REMAINDER(4) => N71, REMAINDER(3) => N70, 
               REMAINDER(2) => N69, REMAINDER(1) => N68, REMAINDER(0) => N67
      );
   lt_94 : process ( X_Logic0_port, VIRTUAL_ADDRESS2_4_port, 
         VIRTUAL_ADDRESS2_3_port, VIRTUAL_ADDRESS2_2_port, 
         VIRTUAL_ADDRESS2_1_port, VIRTUAL_ADDRESS2_0_port, X_Logic1_port )
      variable A : SIGNED( 5 downto 0 );
      variable B : SIGNED( 4 downto 0 );
      variable Z : SIGNED( 0 downto 0 );
   begin
      A := ( X_Logic0_port, VIRTUAL_ADDRESS2_4_port, VIRTUAL_ADDRESS2_3_port, 
            VIRTUAL_ADDRESS2_2_port, VIRTUAL_ADDRESS2_1_port, 
            VIRTUAL_ADDRESS2_0_port );
      B := ( X_Logic0_port, X_Logic1_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port );
      if ( A < B ) then
         Z := ( others => '1' );
      else
         Z := ( others => '0' );
      end if;
      ( 0 => N73 ) <= Z;
   end process;
   
   mod_100 : MOD_UNS_OP
      generic map ( A_width => 6, B_width => 31, REMAINDER_width => 31 )
      port map(
         -- Connections to port 'A'
         A(5) => N92, A(4) => N91, A(3) => N90, A(2) => N89, A(1) => N88, A(0) 
               => N87, 
         -- Connections to port 'B'
         B(30) => X_Logic0_port, B(29) => X_Logic0_port, B(28) => X_Logic0_port
               , B(27) => X_Logic0_port, B(26) => X_Logic0_port, B(25) => 
               X_Logic0_port, B(24) => X_Logic0_port, B(23) => X_Logic0_port, 
               B(22) => X_Logic0_port, B(21) => X_Logic0_port, B(20) => 
               X_Logic0_port, B(19) => X_Logic0_port, B(18) => X_Logic0_port, 
               B(17) => X_Logic0_port, B(16) => X_Logic0_port, B(15) => 
               X_Logic0_port, B(14) => X_Logic0_port, B(13) => X_Logic0_port, 
               B(12) => X_Logic0_port, B(11) => X_Logic0_port, B(10) => 
               X_Logic0_port, B(9) => X_Logic0_port, B(8) => X_Logic0_port, 
               B(7) => X_Logic0_port, B(6) => X_Logic0_port, B(5) => 
               X_Logic1_port, B(4) => X_Logic1_port, B(3) => X_Logic1_port, 
               B(2) => X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
               X_Logic0_port, 
         -- Connections to port 'REMAINDER'
         REMAINDER(30) => n_3163, REMAINDER(29) => n_3164, REMAINDER(28) => 
               n_3165, REMAINDER(27) => n_3166, REMAINDER(26) => n_3167, 
               REMAINDER(25) => n_3168, REMAINDER(24) => n_3169, REMAINDER(23) 
               => n_3170, REMAINDER(22) => n_3171, REMAINDER(21) => n_3172, 
               REMAINDER(20) => n_3173, REMAINDER(19) => n_3174, REMAINDER(18) 
               => n_3175, REMAINDER(17) => n_3176, REMAINDER(16) => n_3177, 
               REMAINDER(15) => n_3178, REMAINDER(14) => n_3179, REMAINDER(13) 
               => n_3180, REMAINDER(12) => n_3181, REMAINDER(11) => n_3182, 
               REMAINDER(10) => n_3183, REMAINDER(9) => n_3184, REMAINDER(8) =>
               n_3185, REMAINDER(7) => n_3186, REMAINDER(6) => n_3187, 
               REMAINDER(5) => N98, REMAINDER(4) => N97, REMAINDER(3) => N96, 
               REMAINDER(2) => N95, REMAINDER(1) => N94, REMAINDER(0) => N93
      );
   lt_103 : process ( X_Logic0_port, VIRTUAL_ADDRESS3_4_port, 
         VIRTUAL_ADDRESS3_3_port, VIRTUAL_ADDRESS3_2_port, 
         VIRTUAL_ADDRESS3_1_port, VIRTUAL_ADDRESS3_0_port, X_Logic1_port )
      variable A : SIGNED( 5 downto 0 );
      variable B : SIGNED( 4 downto 0 );
      variable Z : SIGNED( 0 downto 0 );
   begin
      A := ( X_Logic0_port, VIRTUAL_ADDRESS3_4_port, VIRTUAL_ADDRESS3_3_port, 
            VIRTUAL_ADDRESS3_2_port, VIRTUAL_ADDRESS3_1_port, 
            VIRTUAL_ADDRESS3_0_port );
      B := ( X_Logic0_port, X_Logic1_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port );
      if ( A < B ) then
         Z := ( others => '1' );
      else
         Z := ( others => '0' );
      end if;
      ( 0 => N99 ) <= Z;
   end process;
   
   mod_109 : MOD_UNS_OP
      generic map ( A_width => 6, B_width => 31, REMAINDER_width => 31 )
      port map(
         -- Connections to port 'A'
         A(5) => N118, A(4) => N117, A(3) => N116, A(2) => N115, A(1) => N114, 
               A(0) => N113, 
         -- Connections to port 'B'
         B(30) => X_Logic0_port, B(29) => X_Logic0_port, B(28) => X_Logic0_port
               , B(27) => X_Logic0_port, B(26) => X_Logic0_port, B(25) => 
               X_Logic0_port, B(24) => X_Logic0_port, B(23) => X_Logic0_port, 
               B(22) => X_Logic0_port, B(21) => X_Logic0_port, B(20) => 
               X_Logic0_port, B(19) => X_Logic0_port, B(18) => X_Logic0_port, 
               B(17) => X_Logic0_port, B(16) => X_Logic0_port, B(15) => 
               X_Logic0_port, B(14) => X_Logic0_port, B(13) => X_Logic0_port, 
               B(12) => X_Logic0_port, B(11) => X_Logic0_port, B(10) => 
               X_Logic0_port, B(9) => X_Logic0_port, B(8) => X_Logic0_port, 
               B(7) => X_Logic0_port, B(6) => X_Logic0_port, B(5) => 
               X_Logic1_port, B(4) => X_Logic1_port, B(3) => X_Logic1_port, 
               B(2) => X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
               X_Logic0_port, 
         -- Connections to port 'REMAINDER'
         REMAINDER(30) => n_3188, REMAINDER(29) => n_3189, REMAINDER(28) => 
               n_3190, REMAINDER(27) => n_3191, REMAINDER(26) => n_3192, 
               REMAINDER(25) => n_3193, REMAINDER(24) => n_3194, REMAINDER(23) 
               => n_3195, REMAINDER(22) => n_3196, REMAINDER(21) => n_3197, 
               REMAINDER(20) => n_3198, REMAINDER(19) => n_3199, REMAINDER(18) 
               => n_3200, REMAINDER(17) => n_3201, REMAINDER(16) => n_3202, 
               REMAINDER(15) => n_3203, REMAINDER(14) => n_3204, REMAINDER(13) 
               => n_3205, REMAINDER(12) => n_3206, REMAINDER(11) => n_3207, 
               REMAINDER(10) => n_3208, REMAINDER(9) => n_3209, REMAINDER(8) =>
               n_3210, REMAINDER(7) => n_3211, REMAINDER(6) => n_3212, 
               REMAINDER(5) => N124, REMAINDER(4) => N123, REMAINDER(3) => N122
               , REMAINDER(2) => N121, REMAINDER(1) => N120, REMAINDER(0) => 
               N119
      );
   C570 : GTECH_AND2 port map( A => N125, B => N126, Z => N128);
   C571 : GTECH_AND2 port map( A => N128, B => N127, Z => N129);
   C573 : GTECH_OR2 port map( A => curr_state_2_port, B => curr_state_1_port, Z
                           => N130);
   C574 : GTECH_OR2 port map( A => N130, B => N127, Z => N131);
   C577 : GTECH_OR2 port map( A => curr_state_2_port, B => N126, Z => N133);
   C578 : GTECH_OR2 port map( A => N133, B => curr_state_0_port, Z => N134);
   C582 : GTECH_OR2 port map( A => curr_state_2_port, B => N126, Z => N136);
   C583 : GTECH_OR2 port map( A => N136, B => N127, Z => N137);
   C586 : GTECH_OR2 port map( A => N125, B => curr_state_1_port, Z => N139);
   C587 : GTECH_OR2 port map( A => N139, B => curr_state_0_port, Z => N140);
   ne_153 : process ( N265, N266, N267, N268, N269, N270, N271, N280, N281, 
         N282, N283, N284, N285, N286 )
      variable A : UNSIGNED( 6 downto 0 );
      variable B : UNSIGNED( 6 downto 0 );
      variable Z : UNSIGNED( 0 downto 0 );
   begin
      A := ( N265, N266, N267, N268, N269, N270, N271 );
      B := ( N280, N281, N282, N283, N284, N285, N286 );
      if ( A /= B ) then
         Z := ( others => '1' );
      else
         Z := ( others => '0' );
      end if;
      ( 0 => N147 ) <= Z;
   end process;
   
   eq_156 : process ( N265, N266, N267, N268, N269, N270, N271, N280, N281, 
         N282, N283, N284, N285, N286 )
      variable A : UNSIGNED( 6 downto 0 );
      variable B : UNSIGNED( 6 downto 0 );
      variable Z : UNSIGNED( 0 downto 0 );
   begin
      A := ( N265, N266, N267, N268, N269, N270, N271 );
      B := ( N280, N281, N282, N283, N284, N285, N286 );
      if ( A = B ) then
         Z := ( others => '1' );
      else
         Z := ( others => '0' );
      end if;
      ( 0 => N152 ) <= Z;
   end process;
   
   mod_159 : MOD_UNS_OP
      generic map ( A_width => 7, B_width => 31, REMAINDER_width => 31 )
      port map(
         -- Connections to port 'A'
         A(6) => N159, A(5) => N158, A(4) => N157, A(3) => N156, A(2) => N155, 
               A(1) => N154, A(0) => N153, 
         -- Connections to port 'B'
         B(30) => X_Logic0_port, B(29) => X_Logic0_port, B(28) => X_Logic0_port
               , B(27) => X_Logic0_port, B(26) => X_Logic0_port, B(25) => 
               X_Logic0_port, B(24) => X_Logic0_port, B(23) => X_Logic0_port, 
               B(22) => X_Logic0_port, B(21) => X_Logic0_port, B(20) => 
               X_Logic0_port, B(19) => X_Logic0_port, B(18) => X_Logic0_port, 
               B(17) => X_Logic0_port, B(16) => X_Logic0_port, B(15) => 
               X_Logic0_port, B(14) => X_Logic0_port, B(13) => X_Logic0_port, 
               B(12) => X_Logic0_port, B(11) => X_Logic0_port, B(10) => 
               X_Logic0_port, B(9) => X_Logic0_port, B(8) => X_Logic0_port, 
               B(7) => X_Logic0_port, B(6) => X_Logic0_port, B(5) => 
               X_Logic1_port, B(4) => X_Logic1_port, B(3) => X_Logic1_port, 
               B(2) => X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
               X_Logic0_port, 
         -- Connections to port 'REMAINDER'
         REMAINDER(30) => n_3213, REMAINDER(29) => n_3214, REMAINDER(28) => 
               n_3215, REMAINDER(27) => n_3216, REMAINDER(26) => n_3217, 
               REMAINDER(25) => n_3218, REMAINDER(24) => n_3219, REMAINDER(23) 
               => n_3220, REMAINDER(22) => n_3221, REMAINDER(21) => n_3222, 
               REMAINDER(20) => n_3223, REMAINDER(19) => n_3224, REMAINDER(18) 
               => n_3225, REMAINDER(17) => n_3226, REMAINDER(16) => n_3227, 
               REMAINDER(15) => n_3228, REMAINDER(14) => n_3229, REMAINDER(13) 
               => n_3230, REMAINDER(12) => n_3231, REMAINDER(11) => n_3232, 
               REMAINDER(10) => n_3233, REMAINDER(9) => n_3234, REMAINDER(8) =>
               n_3235, REMAINDER(7) => n_3236, REMAINDER(6) => N166, 
               REMAINDER(5) => N165, REMAINDER(4) => N164, REMAINDER(3) => N163
               , REMAINDER(2) => N162, REMAINDER(1) => N161, REMAINDER(0) => 
               N160
      );
   mod_162 : MOD_UNS_OP
      generic map ( A_width => 7, B_width => 31, REMAINDER_width => 31 )
      port map(
         -- Connections to port 'A'
         A(6) => N176, A(5) => N175, A(4) => N174, A(3) => N173, A(2) => N172, 
               A(1) => N171, A(0) => N170, 
         -- Connections to port 'B'
         B(30) => X_Logic0_port, B(29) => X_Logic0_port, B(28) => X_Logic0_port
               , B(27) => X_Logic0_port, B(26) => X_Logic0_port, B(25) => 
               X_Logic0_port, B(24) => X_Logic0_port, B(23) => X_Logic0_port, 
               B(22) => X_Logic0_port, B(21) => X_Logic0_port, B(20) => 
               X_Logic0_port, B(19) => X_Logic0_port, B(18) => X_Logic0_port, 
               B(17) => X_Logic0_port, B(16) => X_Logic0_port, B(15) => 
               X_Logic0_port, B(14) => X_Logic0_port, B(13) => X_Logic0_port, 
               B(12) => X_Logic0_port, B(11) => X_Logic0_port, B(10) => 
               X_Logic0_port, B(9) => X_Logic0_port, B(8) => X_Logic0_port, 
               B(7) => X_Logic0_port, B(6) => X_Logic0_port, B(5) => 
               X_Logic1_port, B(4) => X_Logic1_port, B(3) => X_Logic1_port, 
               B(2) => X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
               X_Logic0_port, 
         -- Connections to port 'REMAINDER'
         REMAINDER(30) => n_3237, REMAINDER(29) => n_3238, REMAINDER(28) => 
               n_3239, REMAINDER(27) => n_3240, REMAINDER(26) => n_3241, 
               REMAINDER(25) => n_3242, REMAINDER(24) => n_3243, REMAINDER(23) 
               => n_3244, REMAINDER(22) => n_3245, REMAINDER(21) => n_3246, 
               REMAINDER(20) => n_3247, REMAINDER(19) => n_3248, REMAINDER(18) 
               => n_3249, REMAINDER(17) => n_3250, REMAINDER(16) => n_3251, 
               REMAINDER(15) => n_3252, REMAINDER(14) => n_3253, REMAINDER(13) 
               => n_3254, REMAINDER(12) => n_3255, REMAINDER(11) => n_3256, 
               REMAINDER(10) => n_3257, REMAINDER(9) => n_3258, REMAINDER(8) =>
               n_3259, REMAINDER(7) => n_3260, REMAINDER(6) => N183, 
               REMAINDER(5) => N182, REMAINDER(4) => N181, REMAINDER(3) => N180
               , REMAINDER(2) => N179, REMAINDER(1) => N178, REMAINDER(0) => 
               N177
      );
   mod_163 : MOD_UNS_OP
      generic map ( A_width => 7, B_width => 31, REMAINDER_width => 31 )
      port map(
         -- Connections to port 'A'
         A(6) => N190, A(5) => N189, A(4) => N188, A(3) => N187, A(2) => N186, 
               A(1) => N185, A(0) => N184, 
         -- Connections to port 'B'
         B(30) => X_Logic0_port, B(29) => X_Logic0_port, B(28) => X_Logic0_port
               , B(27) => X_Logic0_port, B(26) => X_Logic0_port, B(25) => 
               X_Logic0_port, B(24) => X_Logic0_port, B(23) => X_Logic0_port, 
               B(22) => X_Logic0_port, B(21) => X_Logic0_port, B(20) => 
               X_Logic0_port, B(19) => X_Logic0_port, B(18) => X_Logic0_port, 
               B(17) => X_Logic0_port, B(16) => X_Logic0_port, B(15) => 
               X_Logic0_port, B(14) => X_Logic0_port, B(13) => X_Logic0_port, 
               B(12) => X_Logic0_port, B(11) => X_Logic0_port, B(10) => 
               X_Logic0_port, B(9) => X_Logic0_port, B(8) => X_Logic0_port, 
               B(7) => X_Logic0_port, B(6) => X_Logic0_port, B(5) => 
               X_Logic1_port, B(4) => X_Logic1_port, B(3) => X_Logic1_port, 
               B(2) => X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
               X_Logic0_port, 
         -- Connections to port 'REMAINDER'
         REMAINDER(30) => n_3261, REMAINDER(29) => n_3262, REMAINDER(28) => 
               n_3263, REMAINDER(27) => n_3264, REMAINDER(26) => n_3265, 
               REMAINDER(25) => n_3266, REMAINDER(24) => n_3267, REMAINDER(23) 
               => n_3268, REMAINDER(22) => n_3269, REMAINDER(21) => n_3270, 
               REMAINDER(20) => n_3271, REMAINDER(19) => n_3272, REMAINDER(18) 
               => n_3273, REMAINDER(17) => n_3274, REMAINDER(16) => n_3275, 
               REMAINDER(15) => n_3276, REMAINDER(14) => n_3277, REMAINDER(13) 
               => n_3278, REMAINDER(12) => n_3279, REMAINDER(11) => n_3280, 
               REMAINDER(10) => n_3281, REMAINDER(9) => n_3282, REMAINDER(8) =>
               n_3283, REMAINDER(7) => n_3284, REMAINDER(6) => N197, 
               REMAINDER(5) => N196, REMAINDER(4) => N195, REMAINDER(3) => N194
               , REMAINDER(2) => N193, REMAINDER(1) => N192, REMAINDER(0) => 
               N191
      );
   gt_139 : process ( curr_CANSAVE_1_port, curr_CANSAVE_0_port, X_Logic0_port )
      variable A : UNSIGNED( 1 downto 0 );
      variable B : UNSIGNED( 1 downto 0 );
      variable Z : UNSIGNED( 0 downto 0 );
   begin
      A := ( curr_CANSAVE_1_port, curr_CANSAVE_0_port );
      B := ( X_Logic0_port, X_Logic0_port );
      if ( A > B ) then
         Z := ( others => '1' );
      else
         Z := ( others => '0' );
      end if;
      ( 0 => N200 ) <= Z;
   end process;
   
   mod_147 : MOD_UNS_OP
      generic map ( A_width => 7, B_width => 31, REMAINDER_width => 31 )
      port map(
         -- Connections to port 'A'
         A(6) => N210, A(5) => N209, A(4) => N208, A(3) => N207, A(2) => N206, 
               A(1) => N205, A(0) => N204, 
         -- Connections to port 'B'
         B(30) => X_Logic0_port, B(29) => X_Logic0_port, B(28) => X_Logic0_port
               , B(27) => X_Logic0_port, B(26) => X_Logic0_port, B(25) => 
               X_Logic0_port, B(24) => X_Logic0_port, B(23) => X_Logic0_port, 
               B(22) => X_Logic0_port, B(21) => X_Logic0_port, B(20) => 
               X_Logic0_port, B(19) => X_Logic0_port, B(18) => X_Logic0_port, 
               B(17) => X_Logic0_port, B(16) => X_Logic0_port, B(15) => 
               X_Logic0_port, B(14) => X_Logic0_port, B(13) => X_Logic0_port, 
               B(12) => X_Logic0_port, B(11) => X_Logic0_port, B(10) => 
               X_Logic0_port, B(9) => X_Logic0_port, B(8) => X_Logic0_port, 
               B(7) => X_Logic0_port, B(6) => X_Logic0_port, B(5) => 
               X_Logic1_port, B(4) => X_Logic1_port, B(3) => X_Logic1_port, 
               B(2) => X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
               X_Logic0_port, 
         -- Connections to port 'REMAINDER'
         REMAINDER(30) => n_3285, REMAINDER(29) => n_3286, REMAINDER(28) => 
               n_3287, REMAINDER(27) => n_3288, REMAINDER(26) => n_3289, 
               REMAINDER(25) => n_3290, REMAINDER(24) => n_3291, REMAINDER(23) 
               => n_3292, REMAINDER(22) => n_3293, REMAINDER(21) => n_3294, 
               REMAINDER(20) => n_3295, REMAINDER(19) => n_3296, REMAINDER(18) 
               => n_3297, REMAINDER(17) => n_3298, REMAINDER(16) => n_3299, 
               REMAINDER(15) => n_3300, REMAINDER(14) => n_3301, REMAINDER(13) 
               => n_3302, REMAINDER(12) => n_3303, REMAINDER(11) => n_3304, 
               REMAINDER(10) => n_3305, REMAINDER(9) => n_3306, REMAINDER(8) =>
               n_3307, REMAINDER(7) => n_3308, REMAINDER(6) => N217, 
               REMAINDER(5) => N216, REMAINDER(4) => N215, REMAINDER(3) => N214
               , REMAINDER(2) => N213, REMAINDER(1) => N212, REMAINDER(0) => 
               N211
      );
   mod_150 : MOD_UNS_OP
      generic map ( A_width => 7, B_width => 31, REMAINDER_width => 31 )
      port map(
         -- Connections to port 'A'
         A(6) => N225, A(5) => N224, A(4) => N223, A(3) => N222, A(2) => N221, 
               A(1) => N220, A(0) => N219, 
         -- Connections to port 'B'
         B(30) => X_Logic0_port, B(29) => X_Logic0_port, B(28) => X_Logic0_port
               , B(27) => X_Logic0_port, B(26) => X_Logic0_port, B(25) => 
               X_Logic0_port, B(24) => X_Logic0_port, B(23) => X_Logic0_port, 
               B(22) => X_Logic0_port, B(21) => X_Logic0_port, B(20) => 
               X_Logic0_port, B(19) => X_Logic0_port, B(18) => X_Logic0_port, 
               B(17) => X_Logic0_port, B(16) => X_Logic0_port, B(15) => 
               X_Logic0_port, B(14) => X_Logic0_port, B(13) => X_Logic0_port, 
               B(12) => X_Logic0_port, B(11) => X_Logic0_port, B(10) => 
               X_Logic0_port, B(9) => X_Logic0_port, B(8) => X_Logic0_port, 
               B(7) => X_Logic0_port, B(6) => X_Logic0_port, B(5) => 
               X_Logic1_port, B(4) => X_Logic1_port, B(3) => X_Logic1_port, 
               B(2) => X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
               X_Logic0_port, 
         -- Connections to port 'REMAINDER'
         REMAINDER(30) => n_3309, REMAINDER(29) => n_3310, REMAINDER(28) => 
               n_3311, REMAINDER(27) => n_3312, REMAINDER(26) => n_3313, 
               REMAINDER(25) => n_3314, REMAINDER(24) => n_3315, REMAINDER(23) 
               => n_3316, REMAINDER(22) => n_3317, REMAINDER(21) => n_3318, 
               REMAINDER(20) => n_3319, REMAINDER(19) => n_3320, REMAINDER(18) 
               => n_3321, REMAINDER(17) => n_3322, REMAINDER(16) => n_3323, 
               REMAINDER(15) => n_3324, REMAINDER(14) => n_3325, REMAINDER(13) 
               => n_3326, REMAINDER(12) => n_3327, REMAINDER(11) => n_3328, 
               REMAINDER(10) => n_3329, REMAINDER(9) => n_3330, REMAINDER(8) =>
               n_3331, REMAINDER(7) => n_3332, REMAINDER(6) => N232, 
               REMAINDER(5) => N231, REMAINDER(4) => N230, REMAINDER(3) => N229
               , REMAINDER(2) => N228, REMAINDER(1) => N227, REMAINDER(0) => 
               N226
      );
   next_CANSAVE_reg_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               N260, data_in => N262, synch_clear => X_Logic0_port, 
               synch_preset => X_Logic0_port, synch_toggle => X_Logic0_port, 
               synch_enable => X_Logic0_port, next_state => X_Logic0_port, 
               clocked_on => X_Logic0_port, Q => next_CANSAVE_1_port, QN => 
               n_3333);
   next_CANSAVE_reg_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               N260, data_in => N261, synch_clear => X_Logic0_port, 
               synch_preset => X_Logic0_port, synch_toggle => X_Logic0_port, 
               synch_enable => X_Logic0_port, next_state => X_Logic0_port, 
               clocked_on => X_Logic0_port, Q => next_CANSAVE_0_port, QN => 
               n_3334);
   next_state_reg_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               N233, data_in => N236, synch_clear => X_Logic0_port, 
               synch_preset => X_Logic0_port, synch_toggle => X_Logic0_port, 
               synch_enable => X_Logic0_port, next_state => X_Logic0_port, 
               clocked_on => X_Logic0_port, Q => next_state_2_port, QN => 
               n_3335);
   next_state_reg_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               N233, data_in => N235, synch_clear => X_Logic0_port, 
               synch_preset => X_Logic0_port, synch_toggle => X_Logic0_port, 
               synch_enable => X_Logic0_port, next_state => X_Logic0_port, 
               clocked_on => X_Logic0_port, Q => next_state_1_port, QN => 
               n_3336);
   next_state_reg_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               N233, data_in => N234, synch_clear => X_Logic0_port, 
               synch_preset => X_Logic0_port, synch_toggle => X_Logic0_port, 
               synch_enable => X_Logic0_port, next_state => X_Logic0_port, 
               clocked_on => X_Logic0_port, Q => next_state_0_port, QN => 
               n_3337);
   next_CWP_reg_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               N237, data_in => N244, synch_clear => X_Logic0_port, 
               synch_preset => X_Logic0_port, synch_toggle => X_Logic0_port, 
               synch_enable => X_Logic0_port, next_state => X_Logic0_port, 
               clocked_on => X_Logic0_port, Q => next_CWP_6_port, QN => n_3338
               );
   next_CWP_reg_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               N237, data_in => N243, synch_clear => X_Logic0_port, 
               synch_preset => X_Logic0_port, synch_toggle => X_Logic0_port, 
               synch_enable => X_Logic0_port, next_state => X_Logic0_port, 
               clocked_on => X_Logic0_port, Q => next_CWP_5_port, QN => n_3339
               );
   next_CWP_reg_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               N237, data_in => N242, synch_clear => X_Logic0_port, 
               synch_preset => X_Logic0_port, synch_toggle => X_Logic0_port, 
               synch_enable => X_Logic0_port, next_state => X_Logic0_port, 
               clocked_on => X_Logic0_port, Q => next_CWP_4_port, QN => n_3340
               );
   next_CWP_reg_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               N237, data_in => N241, synch_clear => X_Logic0_port, 
               synch_preset => X_Logic0_port, synch_toggle => X_Logic0_port, 
               synch_enable => X_Logic0_port, next_state => X_Logic0_port, 
               clocked_on => X_Logic0_port, Q => next_CWP_3_port, QN => n_3341
               );
   next_CWP_reg_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               N237, data_in => N240, synch_clear => X_Logic0_port, 
               synch_preset => X_Logic0_port, synch_toggle => X_Logic0_port, 
               synch_enable => X_Logic0_port, next_state => X_Logic0_port, 
               clocked_on => X_Logic0_port, Q => next_CWP_2_port, QN => n_3342
               );
   next_CWP_reg_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               N237, data_in => N239, synch_clear => X_Logic0_port, 
               synch_preset => X_Logic0_port, synch_toggle => X_Logic0_port, 
               synch_enable => X_Logic0_port, next_state => X_Logic0_port, 
               clocked_on => X_Logic0_port, Q => next_CWP_1_port, QN => n_3343
               );
   next_CWP_reg_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               N237, data_in => N238, synch_clear => X_Logic0_port, 
               synch_preset => X_Logic0_port, synch_toggle => X_Logic0_port, 
               synch_enable => X_Logic0_port, next_state => X_Logic0_port, 
               clocked_on => X_Logic0_port, Q => next_CWP_0_port, QN => n_3344
               );
   next_SWP_reg_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               N245, data_in => N252, synch_clear => X_Logic0_port, 
               synch_preset => X_Logic0_port, synch_toggle => X_Logic0_port, 
               synch_enable => X_Logic0_port, next_state => X_Logic0_port, 
               clocked_on => X_Logic0_port, Q => next_SWP_6_port, QN => n_3345
               );
   next_SWP_reg_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               N245, data_in => N251, synch_clear => X_Logic0_port, 
               synch_preset => X_Logic0_port, synch_toggle => X_Logic0_port, 
               synch_enable => X_Logic0_port, next_state => X_Logic0_port, 
               clocked_on => X_Logic0_port, Q => next_SWP_5_port, QN => n_3346
               );
   next_SWP_reg_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               N245, data_in => N250, synch_clear => X_Logic0_port, 
               synch_preset => X_Logic0_port, synch_toggle => X_Logic0_port, 
               synch_enable => X_Logic0_port, next_state => X_Logic0_port, 
               clocked_on => X_Logic0_port, Q => next_SWP_4_port, QN => n_3347
               );
   next_SWP_reg_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               N245, data_in => N249, synch_clear => X_Logic0_port, 
               synch_preset => X_Logic0_port, synch_toggle => X_Logic0_port, 
               synch_enable => X_Logic0_port, next_state => X_Logic0_port, 
               clocked_on => X_Logic0_port, Q => next_SWP_3_port, QN => n_3348
               );
   next_SWP_reg_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               N245, data_in => N248, synch_clear => X_Logic0_port, 
               synch_preset => X_Logic0_port, synch_toggle => X_Logic0_port, 
               synch_enable => X_Logic0_port, next_state => X_Logic0_port, 
               clocked_on => X_Logic0_port, Q => next_SWP_2_port, QN => n_3349
               );
   next_SWP_reg_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               N245, data_in => N247, synch_clear => X_Logic0_port, 
               synch_preset => X_Logic0_port, synch_toggle => X_Logic0_port, 
               synch_enable => X_Logic0_port, next_state => X_Logic0_port, 
               clocked_on => X_Logic0_port, Q => next_SWP_1_port, QN => n_3350
               );
   next_SWP_reg_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               N245, data_in => N246, synch_clear => X_Logic0_port, 
               synch_preset => X_Logic0_port, synch_toggle => X_Logic0_port, 
               synch_enable => X_Logic0_port, next_state => X_Logic0_port, 
               clocked_on => X_Logic0_port, Q => next_SWP_0_port, QN => n_3351
               );
   next_RESTORE_reg_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               N237, data_in => N259, synch_clear => X_Logic0_port, 
               synch_preset => X_Logic0_port, synch_toggle => X_Logic0_port, 
               synch_enable => X_Logic0_port, next_state => X_Logic0_port, 
               clocked_on => X_Logic0_port, Q => next_RESTORE_6_port, QN => 
               n_3352);
   next_RESTORE_reg_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               N237, data_in => N258, synch_clear => X_Logic0_port, 
               synch_preset => X_Logic0_port, synch_toggle => X_Logic0_port, 
               synch_enable => X_Logic0_port, next_state => X_Logic0_port, 
               clocked_on => X_Logic0_port, Q => next_RESTORE_5_port, QN => 
               n_3353);
   next_RESTORE_reg_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               N237, data_in => N257, synch_clear => X_Logic0_port, 
               synch_preset => X_Logic0_port, synch_toggle => X_Logic0_port, 
               synch_enable => X_Logic0_port, next_state => X_Logic0_port, 
               clocked_on => X_Logic0_port, Q => next_RESTORE_4_port, QN => 
               n_3354);
   next_RESTORE_reg_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               N237, data_in => N256, synch_clear => X_Logic0_port, 
               synch_preset => X_Logic0_port, synch_toggle => X_Logic0_port, 
               synch_enable => X_Logic0_port, next_state => X_Logic0_port, 
               clocked_on => X_Logic0_port, Q => next_RESTORE_3_port, QN => 
               n_3355);
   next_RESTORE_reg_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               N237, data_in => N255, synch_clear => X_Logic0_port, 
               synch_preset => X_Logic0_port, synch_toggle => X_Logic0_port, 
               synch_enable => X_Logic0_port, next_state => X_Logic0_port, 
               clocked_on => X_Logic0_port, Q => next_RESTORE_2_port, QN => 
               n_3356);
   next_RESTORE_reg_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               N237, data_in => N254, synch_clear => X_Logic0_port, 
               synch_preset => X_Logic0_port, synch_toggle => X_Logic0_port, 
               synch_enable => X_Logic0_port, next_state => X_Logic0_port, 
               clocked_on => X_Logic0_port, Q => next_RESTORE_1_port, QN => 
               n_3357);
   next_RESTORE_reg_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               N237, data_in => N253, synch_clear => X_Logic0_port, 
               synch_preset => X_Logic0_port, synch_toggle => X_Logic0_port, 
               synch_enable => X_Logic0_port, next_state => X_Logic0_port, 
               clocked_on => X_Logic0_port, Q => next_RESTORE_0_port, QN => 
               n_3358);
   add_88 : process ( X_Logic0_port, VIRTUAL_ADDRESS1_4_port, 
         VIRTUAL_ADDRESS1_3_port, VIRTUAL_ADDRESS1_2_port, 
         VIRTUAL_ADDRESS1_1_port, VIRTUAL_ADDRESS1_0_port, X_Logic1_port )
      variable A : SIGNED( 5 downto 0 );
      variable B : SIGNED( 5 downto 0 );
      variable Z : SIGNED( 5 downto 0 );
   begin
      A := ( X_Logic0_port, VIRTUAL_ADDRESS1_4_port, VIRTUAL_ADDRESS1_3_port, 
            VIRTUAL_ADDRESS1_2_port, VIRTUAL_ADDRESS1_1_port, 
            VIRTUAL_ADDRESS1_0_port );
      B := ( X_Logic1_port, X_Logic1_port, X_Logic1_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port );
      Z := A + B;
      ( N54, N53, N52, N51, N50, N49 ) <= Z;
   end process;
   
   add_97 : process ( X_Logic0_port, VIRTUAL_ADDRESS1_4_port, 
         VIRTUAL_ADDRESS1_3_port, VIRTUAL_ADDRESS1_2_port, 
         VIRTUAL_ADDRESS1_1_port, VIRTUAL_ADDRESS1_0_port, X_Logic1_port )
      variable A : SIGNED( 5 downto 0 );
      variable B : SIGNED( 5 downto 0 );
      variable Z : SIGNED( 5 downto 0 );
   begin
      A := ( X_Logic0_port, VIRTUAL_ADDRESS1_4_port, VIRTUAL_ADDRESS1_3_port, 
            VIRTUAL_ADDRESS1_2_port, VIRTUAL_ADDRESS1_1_port, 
            VIRTUAL_ADDRESS1_0_port );
      B := ( X_Logic1_port, X_Logic1_port, X_Logic1_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port );
      Z := A + B;
      ( N80, N79, N78, N77, N76, N75 ) <= Z;
   end process;
   
   add_106 : process ( X_Logic0_port, VIRTUAL_ADDRESS1_4_port, 
         VIRTUAL_ADDRESS1_3_port, VIRTUAL_ADDRESS1_2_port, 
         VIRTUAL_ADDRESS1_1_port, VIRTUAL_ADDRESS1_0_port, X_Logic1_port )
      variable A : SIGNED( 5 downto 0 );
      variable B : SIGNED( 5 downto 0 );
      variable Z : SIGNED( 5 downto 0 );
   begin
      A := ( X_Logic0_port, VIRTUAL_ADDRESS1_4_port, VIRTUAL_ADDRESS1_3_port, 
            VIRTUAL_ADDRESS1_2_port, VIRTUAL_ADDRESS1_1_port, 
            VIRTUAL_ADDRESS1_0_port );
      B := ( X_Logic1_port, X_Logic1_port, X_Logic1_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port );
      Z := A + B;
      ( N106, N105, N104, N103, N102, N101 ) <= Z;
   end process;
   
   add_91 : process ( VIRTUAL_ADDRESS1_4_port, VIRTUAL_ADDRESS1_3_port, 
         VIRTUAL_ADDRESS1_2_port, VIRTUAL_ADDRESS1_1_port, 
         VIRTUAL_ADDRESS1_0_port, N273, N274, N275, N276, N277, N278 )
      variable A : UNSIGNED( 5 downto 0 );
      variable B : UNSIGNED( 5 downto 0 );
      variable Z : UNSIGNED( 5 downto 0 );
   begin
      A := ( '0', VIRTUAL_ADDRESS1_4_port, VIRTUAL_ADDRESS1_3_port, 
            VIRTUAL_ADDRESS1_2_port, VIRTUAL_ADDRESS1_1_port, 
            VIRTUAL_ADDRESS1_0_port );
      B := ( N273, N274, N275, N276, N277, N278 );
      Z := A + B;
      ( N60, N59, N58, N57, N56, N55 ) <= Z;
   end process;
   
   add_100 : process ( VIRTUAL_ADDRESS2_4_port, VIRTUAL_ADDRESS2_3_port, 
         VIRTUAL_ADDRESS2_2_port, VIRTUAL_ADDRESS2_1_port, 
         VIRTUAL_ADDRESS2_0_port, N273, N274, N275, N276, N277, N278 )
      variable A : UNSIGNED( 5 downto 0 );
      variable B : UNSIGNED( 5 downto 0 );
      variable Z : UNSIGNED( 5 downto 0 );
   begin
      A := ( '0', VIRTUAL_ADDRESS2_4_port, VIRTUAL_ADDRESS2_3_port, 
            VIRTUAL_ADDRESS2_2_port, VIRTUAL_ADDRESS2_1_port, 
            VIRTUAL_ADDRESS2_0_port );
      B := ( N273, N274, N275, N276, N277, N278 );
      Z := A + B;
      ( N86, N85, N84, N83, N82, N81 ) <= Z;
   end process;
   
   add_109 : process ( VIRTUAL_ADDRESS3_4_port, VIRTUAL_ADDRESS3_3_port, 
         VIRTUAL_ADDRESS3_2_port, VIRTUAL_ADDRESS3_1_port, 
         VIRTUAL_ADDRESS3_0_port, N273, N274, N275, N276, N277, N278 )
      variable A : UNSIGNED( 5 downto 0 );
      variable B : UNSIGNED( 5 downto 0 );
      variable Z : UNSIGNED( 5 downto 0 );
   begin
      A := ( '0', VIRTUAL_ADDRESS3_4_port, VIRTUAL_ADDRESS3_3_port, 
            VIRTUAL_ADDRESS3_2_port, VIRTUAL_ADDRESS3_1_port, 
            VIRTUAL_ADDRESS3_0_port );
      B := ( N273, N274, N275, N276, N277, N278 );
      Z := A + B;
      ( N112, N111, N110, N109, N108, N107 ) <= Z;
   end process;
   
   C773 : GTECH_OR3 port map( A => N129, B => N135, C => N141, Z => N237);
   C774 : GTECH_OR2 port map( A => N132, B => N138, Z => N263);
   C815 : GTECH_OR4 port map( A => N129, B => N135, C => N138, D => N141, Z => 
                           N264);
   sub_91 : process ( N60, N59, N58, N57, N56, N55, X_Logic1_port, 
         X_Logic0_port )
      variable A : UNSIGNED( 5 downto 0 );
      variable B : UNSIGNED( 5 downto 0 );
      variable Z : UNSIGNED( 5 downto 0 );
   begin
      A := ( N60, N59, N58, N57, N56, N55 );
      B := ( '0', '0', X_Logic1_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port );
      Z := A - B;
      ( N66, N65, N64, N63, N62, N61 ) <= Z;
   end process;
   
   sub_100 : process ( N86, N85, N84, N83, N82, N81, X_Logic1_port, 
         X_Logic0_port )
      variable A : UNSIGNED( 5 downto 0 );
      variable B : UNSIGNED( 5 downto 0 );
      variable Z : UNSIGNED( 5 downto 0 );
   begin
      A := ( N86, N85, N84, N83, N82, N81 );
      B := ( '0', '0', X_Logic1_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port );
      Z := A - B;
      ( N92, N91, N90, N89, N88, N87 ) <= Z;
   end process;
   
   sub_109 : process ( N112, N111, N110, N109, N108, N107, X_Logic1_port, 
         X_Logic0_port )
      variable A : UNSIGNED( 5 downto 0 );
      variable B : UNSIGNED( 5 downto 0 );
      variable Z : UNSIGNED( 5 downto 0 );
   begin
      A := ( N112, N111, N110, N109, N108, N107 );
      B := ( '0', '0', X_Logic1_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port );
      Z := A - B;
      ( N118, N117, N116, N115, N114, N113 ) <= Z;
   end process;
   
   add_150 : process ( N272, N273, N274, N275, N276, N277, N278, X_Logic1_port,
         X_Logic0_port )
      variable A : UNSIGNED( 6 downto 0 );
      variable B : UNSIGNED( 6 downto 0 );
      variable Z : UNSIGNED( 6 downto 0 );
   begin
      A := ( N272, N273, N274, N275, N276, N277, N278 );
      B := ( '0', '0', X_Logic1_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port );
      Z := A + B;
      ( N225, N224, N223, N222, N221, N220, N219 ) <= Z;
   end process;
   
   sub_162_cf : process ( X_Logic1_port, X_Logic0_port, N265, N266, N267, N268,
         N269, N270, N271 )
      variable A : UNSIGNED( 6 downto 0 );
      variable B : UNSIGNED( 6 downto 0 );
      variable Z : UNSIGNED( 6 downto 0 );
   begin
      A := ( '0', X_Logic1_port, X_Logic0_port, X_Logic1_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port );
      B := ( N265, N266, N267, N268, N269, N270, N271 );
      Z := A + B;
      ( N176, N175, N174, N173, N172, N171, N170 ) <= Z;
   end process;
   
   sub_163_cf : process ( X_Logic1_port, X_Logic0_port, N272, N273, N274, N275,
         N276, N277, N278 )
      variable A : UNSIGNED( 6 downto 0 );
      variable B : UNSIGNED( 6 downto 0 );
      variable Z : UNSIGNED( 6 downto 0 );
   begin
      A := ( '0', X_Logic1_port, X_Logic0_port, X_Logic1_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port );
      B := ( N272, N273, N274, N275, N276, N277, N278 );
      Z := A + B;
      ( N190, N189, N188, N187, N186, N185, N184 ) <= Z;
   end process;
   
   add_154 : process ( curr_CANSAVE_1_port, curr_CANSAVE_0_port, X_Logic1_port 
         )
      variable A : UNSIGNED( 1 downto 0 );
      variable B : UNSIGNED( 1 downto 0 );
      variable Z : UNSIGNED( 1 downto 0 );
   begin
      A := ( curr_CANSAVE_1_port, curr_CANSAVE_0_port );
      B := ( '0', X_Logic1_port );
      Z := A + B;
      ( N150, N149 ) <= Z;
   end process;
   
   sub_141 : process ( curr_CANSAVE_1_port, curr_CANSAVE_0_port, X_Logic1_port 
         )
      variable A : UNSIGNED( 1 downto 0 );
      variable B : UNSIGNED( 1 downto 0 );
      variable Z : UNSIGNED( 1 downto 0 );
   begin
      A := ( curr_CANSAVE_1_port, curr_CANSAVE_0_port );
      B := ( '0', X_Logic1_port );
      Z := A - B;
      ( N203, N202 ) <= Z;
   end process;
   
   add_147 : process ( N272, N273, N274, N275, N276, N277, N278, X_Logic1_port,
         X_Logic0_port )
      variable A : UNSIGNED( 6 downto 0 );
      variable B : UNSIGNED( 6 downto 0 );
      variable Z : UNSIGNED( 6 downto 0 );
   begin
      A := ( N272, N273, N274, N275, N276, N277, N278 );
      B := ( '0', '0', '0', X_Logic1_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port );
      Z := A + B;
      ( N210, N209, N208, N207, N206, N205, N204 ) <= Z;
   end process;
   
   C825 : GTECH_OR4 port map( A => N129, B => N132, C => N135, D => N138, Z => 
                           N279);
   sub_159_cf : process ( X_Logic1_port, X_Logic0_port, N280, N281, N282, N283,
         N284, N285, N286 )
      variable A : UNSIGNED( 6 downto 0 );
      variable B : UNSIGNED( 6 downto 0 );
      variable Z : UNSIGNED( 6 downto 0 );
   begin
      A := ( '0', X_Logic1_port, X_Logic0_port, X_Logic1_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port );
      B := ( N280, N281, N282, N283, N284, N285, N286 );
      Z := A + B;
      ( N159, N158, N157, N156, N155, N154, N153 ) <= Z;
   end process;
   
   C827 : GTECH_OR3 port map( A => N135, B => N138, C => N141, Z => N287);
   C831 : GTECH_OR4 port map( A => N129, B => N132, C => N138, D => N141, Z => 
                           N288);
   C833 : GTECH_OR2 port map( A => N129, B => N132, Z => N289);
   C855_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic1_port, 
         -- Connections to port 'DATA2'
         DATA(1) => ENABLE_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N0, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N1, 
         -- Connections to port 'Z'
         Z(0) => N20 );
   B_0 : GTECH_BUF port map( A => RST, Z => N0);
   B_1 : GTECH_BUF port map( A => N19, Z => N1);
   C856_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 3 )
      port map(
         -- Connections to port 'DATA1'
         DATA(2) => X_Logic0_port, DATA(1) => X_Logic0_port, DATA(0) => 
               X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(5) => next_state_2_port, DATA(4) => next_state_1_port, DATA(3) =>
               next_state_0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N0, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N1, 
         -- Connections to port 'Z'
         Z(2) => N23, Z(1) => N22, Z(0) => N21 );
   C857_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 7 )
      port map(
         -- Connections to port 'DATA1'
         DATA(6) => X_Logic0_port, DATA(5) => X_Logic0_port, DATA(4) => 
               X_Logic0_port, DATA(3) => X_Logic0_port, DATA(2) => 
               X_Logic0_port, DATA(1) => X_Logic0_port, DATA(0) => 
               X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(13) => next_CWP_6_port, DATA(12) => next_CWP_5_port, DATA(11) => 
               next_CWP_4_port, DATA(10) => next_CWP_3_port, DATA(9) => 
               next_CWP_2_port, DATA(8) => next_CWP_1_port, DATA(7) => 
               next_CWP_0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N0, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N1, 
         -- Connections to port 'Z'
         Z(6) => N30, Z(5) => N29, Z(4) => N28, Z(3) => N27, Z(2) => N26, Z(1) 
               => N25, Z(0) => N24 );
   C858_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 7 )
      port map(
         -- Connections to port 'DATA1'
         DATA(6) => X_Logic0_port, DATA(5) => X_Logic0_port, DATA(4) => 
               X_Logic0_port, DATA(3) => X_Logic0_port, DATA(2) => 
               X_Logic0_port, DATA(1) => X_Logic0_port, DATA(0) => 
               X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(13) => next_SWP_6_port, DATA(12) => next_SWP_5_port, DATA(11) => 
               next_SWP_4_port, DATA(10) => next_SWP_3_port, DATA(9) => 
               next_SWP_2_port, DATA(8) => next_SWP_1_port, DATA(7) => 
               next_SWP_0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N0, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N1, 
         -- Connections to port 'Z'
         Z(6) => N37, Z(5) => N36, Z(4) => N35, Z(3) => N34, Z(2) => N33, Z(1) 
               => N32, Z(0) => N31 );
   C859_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 7 )
      port map(
         -- Connections to port 'DATA1'
         DATA(6) => X_Logic0_port, DATA(5) => X_Logic0_port, DATA(4) => 
               X_Logic0_port, DATA(3) => X_Logic0_port, DATA(2) => 
               X_Logic0_port, DATA(1) => X_Logic0_port, DATA(0) => 
               X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(13) => next_RESTORE_6_port, DATA(12) => next_RESTORE_5_port, 
               DATA(11) => next_RESTORE_4_port, DATA(10) => next_RESTORE_3_port
               , DATA(9) => next_RESTORE_2_port, DATA(8) => next_RESTORE_1_port
               , DATA(7) => next_RESTORE_0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N0, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N1, 
         -- Connections to port 'Z'
         Z(6) => N44, Z(5) => N43, Z(4) => N42, Z(3) => N41, Z(2) => N40, Z(1) 
               => N39, Z(0) => N38 );
   C860_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 2 )
      port map(
         -- Connections to port 'DATA1'
         DATA(1) => X_Logic1_port, DATA(0) => X_Logic1_port, 
         -- Connections to port 'DATA2'
         DATA(3) => next_CANSAVE_1_port, DATA(2) => next_CANSAVE_0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N0, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N1, 
         -- Connections to port 'Z'
         Z(1) => N46, Z(0) => N45 );
   C861_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 6 )
      port map(
         -- Connections to port 'DATA1'
         DATA(5) => N54, DATA(4) => N53, DATA(3) => N52, DATA(2) => N51, 
               DATA(1) => N50, DATA(0) => N49, 
         -- Connections to port 'DATA2'
         DATA(11) => N72, DATA(10) => N71, DATA(9) => N70, DATA(8) => N69, 
               DATA(7) => N68, DATA(6) => N67, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N2, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N48, 
         -- Connections to port 'Z'
         Z(5) => PHY_ADDRESS1_5_port, Z(4) => PHY_ADDRESS1_4_port, Z(3) => 
               PHY_ADDRESS1_3_port, Z(2) => PHY_ADDRESS1_2_port, Z(1) => 
               PHY_ADDRESS1_1_port, Z(0) => PHY_ADDRESS1_0_port );
   B_2 : GTECH_BUF port map( A => N47, Z => N2);
   C862_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 6 )
      port map(
         -- Connections to port 'DATA1'
         DATA(5) => N80, DATA(4) => N79, DATA(3) => N78, DATA(2) => N77, 
               DATA(1) => N76, DATA(0) => N75, 
         -- Connections to port 'DATA2'
         DATA(11) => N98, DATA(10) => N97, DATA(9) => N96, DATA(8) => N95, 
               DATA(7) => N94, DATA(6) => N93, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N3, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N74, 
         -- Connections to port 'Z'
         Z(5) => PHY_ADDRESS2_5_port, Z(4) => PHY_ADDRESS2_4_port, Z(3) => 
               PHY_ADDRESS2_3_port, Z(2) => PHY_ADDRESS2_2_port, Z(1) => 
               PHY_ADDRESS2_1_port, Z(0) => PHY_ADDRESS2_0_port );
   B_3 : GTECH_BUF port map( A => N73, Z => N3);
   C863_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 6 )
      port map(
         -- Connections to port 'DATA1'
         DATA(5) => N106, DATA(4) => N105, DATA(3) => N104, DATA(2) => N103, 
               DATA(1) => N102, DATA(0) => N101, 
         -- Connections to port 'DATA2'
         DATA(11) => N124, DATA(10) => N123, DATA(9) => N122, DATA(8) => N121, 
               DATA(7) => N120, DATA(6) => N119, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N4, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N100, 
         -- Connections to port 'Z'
         Z(5) => PHY_ADDRESS3_5_port, Z(4) => PHY_ADDRESS3_4_port, Z(3) => 
               PHY_ADDRESS3_3_port, Z(2) => PHY_ADDRESS3_2_port, Z(1) => 
               PHY_ADDRESS3_1_port, Z(0) => PHY_ADDRESS3_0_port );
   B_4 : GTECH_BUF port map( A => N99, Z => N4);
   C864_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 2 )
      port map(
         -- Connections to port 'DATA1'
         DATA(1) => X_Logic0_port, DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(3) => RET_port, DATA(2) => N143, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N5, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N6, 
         -- Connections to port 'Z'
         Z(1) => N145, Z(0) => N144 );
   B_5 : GTECH_BUF port map( A => CALL_port, Z => N5);
   B_6 : GTECH_BUF port map( A => N142, Z => N6);
   C865_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic1_port, 
         -- Connections to port 'DATA2'
         DATA(1) => N152, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N7, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N148, 
         -- Connections to port 'Z'
         Z(0) => N167 );
   B_7 : GTECH_BUF port map( A => N147, Z => N7);
   I_0 : GTECH_NOT port map( A => N147, Z => N168);
   C867_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => N152, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N7, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N148, 
         -- Connections to port 'Z'
         Z(0) => N169 );
   I_1 : GTECH_NOT port map( A => N200, Z => N218);
   C869_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic1_port, 
         -- Connections to port 'DATA2'
         DATA(1) => N167, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N8, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N9, 
         -- Connections to port 'Z'
         Z(0) => N233 );
   B_8 : GTECH_BUF port map( A => N288, Z => N8);
   B_9 : GTECH_BUF port map( A => N135, Z => N9);
   C870_cell : SELECT_OP
      generic map ( num_inputs => 3, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => ENABLE_port, 
         -- Connections to port 'DATA2'
         DATA(1) => N144, 
         -- Connections to port 'DATA3'
         DATA(2) => X_Logic1_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N10, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N11, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N12, 
         -- Connections to port 'Z'
         Z(0) => N234 );
   B_10 : GTECH_BUF port map( A => N129, Z => N10);
   B_11 : GTECH_BUF port map( A => N132, Z => N11);
   B_12 : GTECH_BUF port map( A => N287, Z => N12);
   C871_cell : SELECT_OP
      generic map ( num_inputs => 5, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => N145, 
         -- Connections to port 'DATA3'
         DATA(2) => N168, 
         -- Connections to port 'DATA4'
         DATA(3) => N198, 
         -- Connections to port 'DATA5'
         DATA(4) => N218, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N10, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N11, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N9, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N13, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N14, 
         -- Connections to port 'Z'
         Z(0) => N235 );
   B_13 : GTECH_BUF port map( A => N138, Z => N13);
   B_14 : GTECH_BUF port map( A => N141, Z => N14);
   C872_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => CALL_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N15, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N11, 
         -- Connections to port 'Z'
         Z(0) => N236 );
   B_15 : GTECH_BUF port map( A => N264, Z => N15);
   C873_cell : SELECT_OP
      generic map ( num_inputs => 3, input_width => 7 )
      port map(
         -- Connections to port 'DATA1'
         DATA(6) => X_Logic0_port, DATA(5) => X_Logic0_port, DATA(4) => 
               X_Logic0_port, DATA(3) => X_Logic0_port, DATA(2) => 
               X_Logic0_port, DATA(1) => X_Logic0_port, DATA(0) => 
               X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(13) => N197, DATA(12) => N196, DATA(11) => N195, DATA(10) => N194
               , DATA(9) => N193, DATA(8) => N192, DATA(7) => N191, 
         -- Connections to port 'DATA3'
         DATA(20) => N232, DATA(19) => N231, DATA(18) => N230, DATA(17) => N229
               , DATA(16) => N228, DATA(15) => N227, DATA(14) => N226, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N10, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N9, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N14, 
         -- Connections to port 'Z'
         Z(6) => N244, Z(5) => N243, Z(4) => N242, Z(3) => N241, Z(2) => N240, 
               Z(1) => N239, Z(0) => N238 );
   C874_cell : SELECT_OP
      generic map ( num_inputs => 4, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic1_port, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'DATA3'
         DATA(2) => N169, 
         -- Connections to port 'DATA4'
         DATA(3) => N218, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N10, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N16, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N9, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N14, 
         -- Connections to port 'Z'
         Z(0) => N245 );
   B_16 : GTECH_BUF port map( A => N263, Z => N16);
   C875_cell : SELECT_OP
      generic map ( num_inputs => 3, input_width => 7 )
      port map(
         -- Connections to port 'DATA1'
         DATA(6) => X_Logic0_port, DATA(5) => X_Logic0_port, DATA(4) => 
               X_Logic0_port, DATA(3) => X_Logic0_port, DATA(2) => 
               X_Logic0_port, DATA(1) => X_Logic0_port, DATA(0) => 
               X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(13) => N166, DATA(12) => N165, DATA(11) => N164, DATA(10) => N163
               , DATA(9) => N162, DATA(8) => N161, DATA(7) => N160, 
         -- Connections to port 'DATA3'
         DATA(20) => N217, DATA(19) => N216, DATA(18) => N215, DATA(17) => N214
               , DATA(16) => N213, DATA(15) => N212, DATA(14) => N211, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N10, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N9, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N14, 
         -- Connections to port 'Z'
         Z(6) => N252, Z(5) => N251, Z(4) => N250, Z(3) => N249, Z(2) => N248, 
               Z(1) => N247, Z(0) => N246 );
   C876_cell : SELECT_OP
      generic map ( num_inputs => 3, input_width => 7 )
      port map(
         -- Connections to port 'DATA1'
         DATA(6) => X_Logic0_port, DATA(5) => X_Logic0_port, DATA(4) => 
               X_Logic0_port, DATA(3) => X_Logic0_port, DATA(2) => 
               X_Logic0_port, DATA(1) => X_Logic0_port, DATA(0) => 
               X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(13) => N183, DATA(12) => N182, DATA(11) => N181, DATA(10) => N180
               , DATA(9) => N179, DATA(8) => N178, DATA(7) => N177, 
         -- Connections to port 'DATA3'
         DATA(20) => N272, DATA(19) => N273, DATA(18) => N274, DATA(17) => N275
               , DATA(16) => N276, DATA(15) => N277, DATA(14) => N278, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N10, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N9, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N14, 
         -- Connections to port 'Z'
         Z(6) => N259, Z(5) => N258, Z(4) => N257, Z(3) => N256, Z(2) => N255, 
               Z(1) => N254, Z(0) => N253 );
   C877_cell : SELECT_OP
      generic map ( num_inputs => 4, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic1_port, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'DATA3'
         DATA(2) => N147, 
         -- Connections to port 'DATA4'
         DATA(3) => N200, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N10, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N16, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N9, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N14, 
         -- Connections to port 'Z'
         Z(0) => N260 );
   C878_cell : SELECT_OP
      generic map ( num_inputs => 3, input_width => 2 )
      port map(
         -- Connections to port 'DATA1'
         DATA(1) => X_Logic1_port, DATA(0) => X_Logic1_port, 
         -- Connections to port 'DATA2'
         DATA(3) => N150, DATA(2) => N149, 
         -- Connections to port 'DATA3'
         DATA(5) => N203, DATA(4) => N202, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N10, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N9, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N14, 
         -- Connections to port 'Z'
         Z(1) => N262, Z(0) => N261 );
   C879_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => READ1_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N15, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N11, 
         -- Connections to port 'Z'
         Z(0) => RD1_port );
   C880_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => READ2_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N15, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N11, 
         -- Connections to port 'Z'
         Z(0) => RD2_port );
   C881_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => WRITE_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N15, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N11, 
         -- Connections to port 'Z'
         Z(0) => WR_port );
   C882_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => N169, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N8, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N9, 
         -- Connections to port 'Z'
         Z(0) => FILL_port );
   C883_cell : SELECT_OP
      generic map ( num_inputs => 4, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => N169, 
         -- Connections to port 'DATA3'
         DATA(2) => X_Logic1_port, 
         -- Connections to port 'DATA4'
         DATA(3) => N218, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N17, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N9, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N13, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N14, 
         -- Connections to port 'Z'
         Z(0) => STALL_port );
   B_17 : GTECH_BUF port map( A => N289, Z => N17);
   C884_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => N218, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N18, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N14, 
         -- Connections to port 'Z'
         Z(0) => SPILL_port );
   B_18 : GTECH_BUF port map( A => N279, Z => N18);
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   I_2 : GTECH_NOT port map( A => RST, Z => N19);
   I_3 : GTECH_NOT port map( A => N47, Z => N48);
   B_19 : GTECH_BUF port map( A => N47, Z => net30);
   B_20 : GTECH_BUF port map( A => N48, Z => net31);
   I_4 : GTECH_NOT port map( A => N73, Z => N74);
   B_21 : GTECH_BUF port map( A => N73, Z => net33);
   B_22 : GTECH_BUF port map( A => N74, Z => net34);
   I_5 : GTECH_NOT port map( A => N99, Z => N100);
   B_23 : GTECH_BUF port map( A => N99, Z => net36);
   B_24 : GTECH_BUF port map( A => N100, Z => net37);
   I_6 : GTECH_NOT port map( A => curr_state_2_port, Z => N125);
   I_7 : GTECH_NOT port map( A => curr_state_1_port, Z => N126);
   I_8 : GTECH_NOT port map( A => curr_state_0_port, Z => N127);
   I_9 : GTECH_NOT port map( A => N131, Z => N132);
   I_10 : GTECH_NOT port map( A => N134, Z => N135);
   I_11 : GTECH_NOT port map( A => N137, Z => N138);
   I_12 : GTECH_NOT port map( A => N140, Z => N141);
   I_13 : GTECH_NOT port map( A => CALL_port, Z => N142);
   I_14 : GTECH_NOT port map( A => RET_port, Z => N143);
   B_25 : GTECH_BUF port map( A => N135, Z => N146);
   I_15 : GTECH_NOT port map( A => N147, Z => N148);
   C929 : GTECH_AND2 port map( A => N146, B => N147, Z => n_3359);
   C930 : GTECH_AND2 port map( A => N146, B => N148, Z => N151);
   C932 : GTECH_AND2 port map( A => N151, B => N152, Z => n_3360);
   I_16 : GTECH_NOT port map( A => ACK, Z => N198);
   B_26 : GTECH_BUF port map( A => N141, Z => N199);
   I_17 : GTECH_NOT port map( A => N200, Z => N201);
   C938 : GTECH_AND2 port map( A => N199, B => N200, Z => n_3361);
   C939 : GTECH_AND2 port map( A => N199, B => N201, Z => n_3362);

end SYN_HLSM;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_topLevel_1.all;

entity topLevel_1 is

   port( CALL, RET, CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, 
         ADD_RD1, ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
         std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector (31
         downto 0);  ACK : in std_logic;  SPILL, FILL, STALL : out std_logic);

end topLevel_1;

architecture SYN_STRUCT of topLevel_1 is

   component register_file_WORD_SIZE32_ADDR_SIZE6
      port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
            ADD_RD2 : in std_logic_vector (5 downto 0);  DATAIN : in 
            std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component RMU_M8_N8_F3_VIRTUAL_ADDR_SIZE5_PHY_ADDR_SIZE6
      port( CALL, RET : in std_logic;  STALL : out std_logic;  READ1, READ2, 
            WRITE : in std_logic;  RD1, RD2, WR : out std_logic;  ENABLE, RST, 
            CLK : in std_logic;  SPILL, FILL : out std_logic;  ACK : in 
            std_logic;  PHY_ADDRESS1, PHY_ADDRESS2, PHY_ADDRESS3 : out 
            std_logic_vector (5 downto 0);  VIRTUAL_ADDRESS1, VIRTUAL_ADDRESS2,
            VIRTUAL_ADDRESS3 : in std_logic_vector (4 downto 0));
   end component;
   
   signal BYPASSED_RD1, BYPASSED_RD2, BYPASSED_WR, PHY_ADDRESS1_5_port, 
      PHY_ADDRESS1_4_port, PHY_ADDRESS1_3_port, PHY_ADDRESS1_2_port, 
      PHY_ADDRESS1_1_port, PHY_ADDRESS1_0_port, PHY_ADDRESS2_5_port, 
      PHY_ADDRESS2_4_port, PHY_ADDRESS2_3_port, PHY_ADDRESS2_2_port, 
      PHY_ADDRESS2_1_port, PHY_ADDRESS2_0_port, PHY_ADDRESS3_5_port, 
      PHY_ADDRESS3_4_port, PHY_ADDRESS3_3_port, PHY_ADDRESS3_2_port, 
      PHY_ADDRESS3_1_port, PHY_ADDRESS3_0_port : std_logic;

begin
   
   RegManUn : RMU_M8_N8_F3_VIRTUAL_ADDR_SIZE5_PHY_ADDR_SIZE6 port map( CALL => 
                           CALL, RET => RET, STALL => STALL, READ1 => RD1, 
                           READ2 => RD2, WRITE => WR, RD1 => BYPASSED_RD1, RD2 
                           => BYPASSED_RD2, WR => BYPASSED_WR, ENABLE => ENABLE
                           , RST => RESET, CLK => CLK, SPILL => SPILL, FILL => 
                           FILL, ACK => ACK, PHY_ADDRESS1(5) => 
                           PHY_ADDRESS1_5_port, PHY_ADDRESS1(4) => 
                           PHY_ADDRESS1_4_port, PHY_ADDRESS1(3) => 
                           PHY_ADDRESS1_3_port, PHY_ADDRESS1(2) => 
                           PHY_ADDRESS1_2_port, PHY_ADDRESS1(1) => 
                           PHY_ADDRESS1_1_port, PHY_ADDRESS1(0) => 
                           PHY_ADDRESS1_0_port, PHY_ADDRESS2(5) => 
                           PHY_ADDRESS2_5_port, PHY_ADDRESS2(4) => 
                           PHY_ADDRESS2_4_port, PHY_ADDRESS2(3) => 
                           PHY_ADDRESS2_3_port, PHY_ADDRESS2(2) => 
                           PHY_ADDRESS2_2_port, PHY_ADDRESS2(1) => 
                           PHY_ADDRESS2_1_port, PHY_ADDRESS2(0) => 
                           PHY_ADDRESS2_0_port, PHY_ADDRESS3(5) => 
                           PHY_ADDRESS3_5_port, PHY_ADDRESS3(4) => 
                           PHY_ADDRESS3_4_port, PHY_ADDRESS3(3) => 
                           PHY_ADDRESS3_3_port, PHY_ADDRESS3(2) => 
                           PHY_ADDRESS3_2_port, PHY_ADDRESS3(1) => 
                           PHY_ADDRESS3_1_port, PHY_ADDRESS3(0) => 
                           PHY_ADDRESS3_0_port, VIRTUAL_ADDRESS1(4) => 
                           ADD_WR(4), VIRTUAL_ADDRESS1(3) => ADD_WR(3), 
                           VIRTUAL_ADDRESS1(2) => ADD_WR(2), 
                           VIRTUAL_ADDRESS1(1) => ADD_WR(1), 
                           VIRTUAL_ADDRESS1(0) => ADD_WR(0), 
                           VIRTUAL_ADDRESS2(4) => ADD_RD1(4), 
                           VIRTUAL_ADDRESS2(3) => ADD_RD1(3), 
                           VIRTUAL_ADDRESS2(2) => ADD_RD1(2), 
                           VIRTUAL_ADDRESS2(1) => ADD_RD1(1), 
                           VIRTUAL_ADDRESS2(0) => ADD_RD1(0), 
                           VIRTUAL_ADDRESS3(4) => ADD_RD2(4), 
                           VIRTUAL_ADDRESS3(3) => ADD_RD2(3), 
                           VIRTUAL_ADDRESS3(2) => ADD_RD2(2), 
                           VIRTUAL_ADDRESS3(1) => ADD_RD2(1), 
                           VIRTUAL_ADDRESS3(0) => ADD_RD2(0));
   RegFile : register_file_WORD_SIZE32_ADDR_SIZE6 port map( CLK => CLK, RESET 
                           => RESET, ENABLE => ENABLE, RD1 => BYPASSED_RD1, RD2
                           => BYPASSED_RD2, WR => BYPASSED_WR, ADD_WR(5) => 
                           PHY_ADDRESS1_5_port, ADD_WR(4) => 
                           PHY_ADDRESS1_4_port, ADD_WR(3) => 
                           PHY_ADDRESS1_3_port, ADD_WR(2) => 
                           PHY_ADDRESS1_2_port, ADD_WR(1) => 
                           PHY_ADDRESS1_1_port, ADD_WR(0) => 
                           PHY_ADDRESS1_0_port, ADD_RD1(5) => 
                           PHY_ADDRESS2_5_port, ADD_RD1(4) => 
                           PHY_ADDRESS2_4_port, ADD_RD1(3) => 
                           PHY_ADDRESS2_3_port, ADD_RD1(2) => 
                           PHY_ADDRESS2_2_port, ADD_RD1(1) => 
                           PHY_ADDRESS2_1_port, ADD_RD1(0) => 
                           PHY_ADDRESS2_0_port, ADD_RD2(5) => 
                           PHY_ADDRESS3_5_port, ADD_RD2(4) => 
                           PHY_ADDRESS3_4_port, ADD_RD2(3) => 
                           PHY_ADDRESS3_3_port, ADD_RD2(2) => 
                           PHY_ADDRESS3_2_port, ADD_RD2(1) => 
                           PHY_ADDRESS3_1_port, ADD_RD2(0) => 
                           PHY_ADDRESS3_0_port, DATAIN(31) => DATAIN(31), 
                           DATAIN(30) => DATAIN(30), DATAIN(29) => DATAIN(29), 
                           DATAIN(28) => DATAIN(28), DATAIN(27) => DATAIN(27), 
                           DATAIN(26) => DATAIN(26), DATAIN(25) => DATAIN(25), 
                           DATAIN(24) => DATAIN(24), DATAIN(23) => DATAIN(23), 
                           DATAIN(22) => DATAIN(22), DATAIN(21) => DATAIN(21), 
                           DATAIN(20) => DATAIN(20), DATAIN(19) => DATAIN(19), 
                           DATAIN(18) => DATAIN(18), DATAIN(17) => DATAIN(17), 
                           DATAIN(16) => DATAIN(16), DATAIN(15) => DATAIN(15), 
                           DATAIN(14) => DATAIN(14), DATAIN(13) => DATAIN(13), 
                           DATAIN(12) => DATAIN(12), DATAIN(11) => DATAIN(11), 
                           DATAIN(10) => DATAIN(10), DATAIN(9) => DATAIN(9), 
                           DATAIN(8) => DATAIN(8), DATAIN(7) => DATAIN(7), 
                           DATAIN(6) => DATAIN(6), DATAIN(5) => DATAIN(5), 
                           DATAIN(4) => DATAIN(4), DATAIN(3) => DATAIN(3), 
                           DATAIN(2) => DATAIN(2), DATAIN(1) => DATAIN(1), 
                           DATAIN(0) => DATAIN(0), OUT1(31) => OUT1(31), 
                           OUT1(30) => OUT1(30), OUT1(29) => OUT1(29), OUT1(28)
                           => OUT1(28), OUT1(27) => OUT1(27), OUT1(26) => 
                           OUT1(26), OUT1(25) => OUT1(25), OUT1(24) => OUT1(24)
                           , OUT1(23) => OUT1(23), OUT1(22) => OUT1(22), 
                           OUT1(21) => OUT1(21), OUT1(20) => OUT1(20), OUT1(19)
                           => OUT1(19), OUT1(18) => OUT1(18), OUT1(17) => 
                           OUT1(17), OUT1(16) => OUT1(16), OUT1(15) => OUT1(15)
                           , OUT1(14) => OUT1(14), OUT1(13) => OUT1(13), 
                           OUT1(12) => OUT1(12), OUT1(11) => OUT1(11), OUT1(10)
                           => OUT1(10), OUT1(9) => OUT1(9), OUT1(8) => OUT1(8),
                           OUT1(7) => OUT1(7), OUT1(6) => OUT1(6), OUT1(5) => 
                           OUT1(5), OUT1(4) => OUT1(4), OUT1(3) => OUT1(3), 
                           OUT1(2) => OUT1(2), OUT1(1) => OUT1(1), OUT1(0) => 
                           OUT1(0), OUT2(31) => OUT2(31), OUT2(30) => OUT2(30),
                           OUT2(29) => OUT2(29), OUT2(28) => OUT2(28), OUT2(27)
                           => OUT2(27), OUT2(26) => OUT2(26), OUT2(25) => 
                           OUT2(25), OUT2(24) => OUT2(24), OUT2(23) => OUT2(23)
                           , OUT2(22) => OUT2(22), OUT2(21) => OUT2(21), 
                           OUT2(20) => OUT2(20), OUT2(19) => OUT2(19), OUT2(18)
                           => OUT2(18), OUT2(17) => OUT2(17), OUT2(16) => 
                           OUT2(16), OUT2(15) => OUT2(15), OUT2(14) => OUT2(14)
                           , OUT2(13) => OUT2(13), OUT2(12) => OUT2(12), 
                           OUT2(11) => OUT2(11), OUT2(10) => OUT2(10), OUT2(9) 
                           => OUT2(9), OUT2(8) => OUT2(8), OUT2(7) => OUT2(7), 
                           OUT2(6) => OUT2(6), OUT2(5) => OUT2(5), OUT2(4) => 
                           OUT2(4), OUT2(3) => OUT2(3), OUT2(2) => OUT2(2), 
                           OUT2(1) => OUT2(1), OUT2(0) => OUT2(0));

end SYN_STRUCT;

library IEEE;

use IEEE.std_logic_1164.all;
entity SELECT_OP is
   generic ( num_inputs, input_width : integer );
   port(
      DATA : in std_logic_vector( num_inputs  * input_width - 1 downto 0 );
      CONTROL : in std_logic_vector( num_inputs - 1 downto 0 );
      Z : out std_logic_vector( input_width - 1 downto 0 )
   );
end SELECT_OP;

architecture RTL of SELECT_OP is
begin

   process ( DATA, CONTROL )
      variable index, high, low : integer;
   begin
   
      --  Initialize variables
      index := 0;
      
      -- Loop over the values of the control inputs
      for_loop : for i in CONTROL'range loop
      
         if ( CONTROL(i) = '1' ) then
         
            index := i;
            exit for_loop;
            
         end if;
         
      end loop;
      
      -- Store the corresponding data lines into the output
      low := input_width * index;
      high := low + input_width - 1;
      Z <= DATA( high downto low );
   
   end process;
   
end RTL;

library IEEE;

use IEEE.std_logic_1164.all;

entity SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT is
   generic ( ac_as_q, ac_as_qn, sc_ss_q : integer );
   port(
      clear, preset, enable, data_in, synch_clear, synch_preset, synch_toggle, 
         synch_enable, next_state, clocked_on : in std_logic;
      Q, QN : buffer std_logic
   );
end SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT;

architecture RTL of SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT is
begin

   process ( preset, clear, enable, data_in, clocked_on )
   begin
   
            -- Check the value of inputs (asynchronous first)
            if ( ( ( preset /= '1' ) and ( preset /= '0' ) ) or ( ( clear /= 
                     '1' ) and ( clear /= '0' ) )  ) then
               Q <= 'X';
            elsif ( clear = '1' and preset = '1' ) then
               case ac_as_q is
                  when 2 =>
                     Q <= '1';
                  when 1 =>
                     Q <= '0';
                  when others =>
                     Q <= 'X';
               end case;
               case ac_as_qn is
                  when 2 =>
                     QN <= '1';
                  when 1 =>
                     QN <= '0';
                  when others =>
                     QN <= 'X';
               end case;
            elsif ( clear = '1' ) then
               Q <= '0';
            elsif ( preset = '1' ) then
               Q <= '1';
            elsif ( ( enable /= '1' ) and ( enable /= '0' ) ) then
               Q <= 'X';
            elsif ( enable = '1' ) then
               Q <= data_in;
            elsif ( ( clocked_on /= '1' ) and ( clocked_on /= '0' ) ) then
               Q <= 'X';
            elsif ( clocked_on'event and clocked_on = '1' ) then
         if ( ( ( synch_preset /= '1' ) and ( synch_preset /= '0' ) ) or ( ( 
                  synch_clear /= '1' ) and ( synch_clear /= '0' ) )  ) then
            Q <= 'X';
         elsif ( synch_clear = '1' and synch_preset = '1' ) then
            case sc_ss_q is
               when 2 =>
                  Q <= '1';
               when 1 =>
                  Q <= '0';
               when others =>
                  Q <= 'X';
            end case;
         elsif ( synch_clear = '1' ) then
            Q <= '0';
         elsif ( synch_preset = '1' ) then
            Q <= '1';
         elsif ( ( ( synch_toggle /= '1' ) and ( synch_toggle /= '0' ) ) or ( (
                  synch_enable /= '1' ) and ( synch_enable /= '0' ) )  ) then
            Q <= 'X';
         elsif ( synch_enable = '1' and synch_toggle = '1' ) then
            Q <= 'X';
         elsif ( synch_toggle = '1' ) then
            Q <= QN;
         elsif ( synch_enable = '1' ) then
            Q <= next_state;
         end if;
      end if;
   
   end process;

end RTL;
