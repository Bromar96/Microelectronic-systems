
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_P4Adder is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_P4Adder;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_95 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_95;

architecture SYN_ARCH2 of ND2_95 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_94 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_94;

architecture SYN_ARCH2 of ND2_94 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_93 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_93;

architecture SYN_ARCH2 of ND2_93 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_92 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_92;

architecture SYN_ARCH2 of ND2_92 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_91 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_91;

architecture SYN_ARCH2 of ND2_91 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_90 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_90;

architecture SYN_ARCH2 of ND2_90 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_89 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_89;

architecture SYN_ARCH2 of ND2_89 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_88 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_88;

architecture SYN_ARCH2 of ND2_88 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_87 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_87;

architecture SYN_ARCH2 of ND2_87 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_86 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_86;

architecture SYN_ARCH2 of ND2_86 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_85 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_85;

architecture SYN_ARCH2 of ND2_85 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_84 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_84;

architecture SYN_ARCH2 of ND2_84 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_83 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_83;

architecture SYN_ARCH2 of ND2_83 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_82 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_82;

architecture SYN_ARCH2 of ND2_82 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_81 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_81;

architecture SYN_ARCH2 of ND2_81 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_80 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_80;

architecture SYN_ARCH2 of ND2_80 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_79 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_79;

architecture SYN_ARCH2 of ND2_79 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_78 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_78;

architecture SYN_ARCH2 of ND2_78 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_77 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_77;

architecture SYN_ARCH2 of ND2_77 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_76 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_76;

architecture SYN_ARCH2 of ND2_76 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_75 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_75;

architecture SYN_ARCH2 of ND2_75 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_74 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_74;

architecture SYN_ARCH2 of ND2_74 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_73 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_73;

architecture SYN_ARCH2 of ND2_73 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_72 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_72;

architecture SYN_ARCH2 of ND2_72 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_71 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_71;

architecture SYN_ARCH2 of ND2_71 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_70 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_70;

architecture SYN_ARCH2 of ND2_70 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_69 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_69;

architecture SYN_ARCH2 of ND2_69 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_68 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_68;

architecture SYN_ARCH2 of ND2_68 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_67 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_67;

architecture SYN_ARCH2 of ND2_67 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_66 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_66;

architecture SYN_ARCH2 of ND2_66 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_65 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_65;

architecture SYN_ARCH2 of ND2_65 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_64 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_64;

architecture SYN_ARCH2 of ND2_64 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_63 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_63;

architecture SYN_ARCH2 of ND2_63 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_62 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_62;

architecture SYN_ARCH2 of ND2_62 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_61 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_61;

architecture SYN_ARCH2 of ND2_61 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_60 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_60;

architecture SYN_ARCH2 of ND2_60 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_59 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_59;

architecture SYN_ARCH2 of ND2_59 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_58 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_58;

architecture SYN_ARCH2 of ND2_58 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_57 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_57;

architecture SYN_ARCH2 of ND2_57 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_56 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_56;

architecture SYN_ARCH2 of ND2_56 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_55 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_55;

architecture SYN_ARCH2 of ND2_55 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_54 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_54;

architecture SYN_ARCH2 of ND2_54 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_53 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_53;

architecture SYN_ARCH2 of ND2_53 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_52 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_52;

architecture SYN_ARCH2 of ND2_52 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_51 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_51;

architecture SYN_ARCH2 of ND2_51 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_50 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_50;

architecture SYN_ARCH2 of ND2_50 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_49 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_49;

architecture SYN_ARCH2 of ND2_49 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_48 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_48;

architecture SYN_ARCH2 of ND2_48 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_47 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_47;

architecture SYN_ARCH2 of ND2_47 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_46 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_46;

architecture SYN_ARCH2 of ND2_46 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_45 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_45;

architecture SYN_ARCH2 of ND2_45 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_44 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_44;

architecture SYN_ARCH2 of ND2_44 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_43 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_43;

architecture SYN_ARCH2 of ND2_43 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_42 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_42;

architecture SYN_ARCH2 of ND2_42 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_41 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_41;

architecture SYN_ARCH2 of ND2_41 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_40 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_40;

architecture SYN_ARCH2 of ND2_40 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_39 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_39;

architecture SYN_ARCH2 of ND2_39 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_38 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_38;

architecture SYN_ARCH2 of ND2_38 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_37 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_37;

architecture SYN_ARCH2 of ND2_37 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_36 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_36;

architecture SYN_ARCH2 of ND2_36 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_35 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_35;

architecture SYN_ARCH2 of ND2_35 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_34 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_34;

architecture SYN_ARCH2 of ND2_34 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_33 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_33;

architecture SYN_ARCH2 of ND2_33 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_32 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_32;

architecture SYN_ARCH2 of ND2_32 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_31 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_31;

architecture SYN_ARCH2 of ND2_31 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_30 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_30;

architecture SYN_ARCH2 of ND2_30 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_29 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_29;

architecture SYN_ARCH2 of ND2_29 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_28 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_28;

architecture SYN_ARCH2 of ND2_28 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_27 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_27;

architecture SYN_ARCH2 of ND2_27 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_26 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_26;

architecture SYN_ARCH2 of ND2_26 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_25 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_25;

architecture SYN_ARCH2 of ND2_25 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_24 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_24;

architecture SYN_ARCH2 of ND2_24 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_23 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_23;

architecture SYN_ARCH2 of ND2_23 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_22 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_22;

architecture SYN_ARCH2 of ND2_22 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_21 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_21;

architecture SYN_ARCH2 of ND2_21 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_20 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_20;

architecture SYN_ARCH2 of ND2_20 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_19 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_19;

architecture SYN_ARCH2 of ND2_19 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_18 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_18;

architecture SYN_ARCH2 of ND2_18 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_17 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_17;

architecture SYN_ARCH2 of ND2_17 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_16 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_16;

architecture SYN_ARCH2 of ND2_16 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_15 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_15;

architecture SYN_ARCH2 of ND2_15 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_14 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_14;

architecture SYN_ARCH2 of ND2_14 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_13 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_13;

architecture SYN_ARCH2 of ND2_13 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_12 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_12;

architecture SYN_ARCH2 of ND2_12 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_11 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_11;

architecture SYN_ARCH2 of ND2_11 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_10 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_10;

architecture SYN_ARCH2 of ND2_10 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_9 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_9;

architecture SYN_ARCH2 of ND2_9 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_8 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_8;

architecture SYN_ARCH2 of ND2_8 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_7 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_7;

architecture SYN_ARCH2 of ND2_7 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_6 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_6;

architecture SYN_ARCH2 of ND2_6 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_5 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_5;

architecture SYN_ARCH2 of ND2_5 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_4 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_4;

architecture SYN_ARCH2 of ND2_4 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_3 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_3;

architecture SYN_ARCH2 of ND2_3 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_2 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_2;

architecture SYN_ARCH2 of ND2_2 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_1 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_1;

architecture SYN_ARCH2 of ND2_1 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity IV_31 is

   port( A : in std_logic;  Y : out std_logic);

end IV_31;

architecture SYN_BEHAVIORAL of IV_31 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity IV_30 is

   port( A : in std_logic;  Y : out std_logic);

end IV_30;

architecture SYN_BEHAVIORAL of IV_30 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity IV_29 is

   port( A : in std_logic;  Y : out std_logic);

end IV_29;

architecture SYN_BEHAVIORAL of IV_29 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity IV_28 is

   port( A : in std_logic;  Y : out std_logic);

end IV_28;

architecture SYN_BEHAVIORAL of IV_28 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity IV_27 is

   port( A : in std_logic;  Y : out std_logic);

end IV_27;

architecture SYN_BEHAVIORAL of IV_27 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity IV_26 is

   port( A : in std_logic;  Y : out std_logic);

end IV_26;

architecture SYN_BEHAVIORAL of IV_26 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity IV_25 is

   port( A : in std_logic;  Y : out std_logic);

end IV_25;

architecture SYN_BEHAVIORAL of IV_25 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity IV_24 is

   port( A : in std_logic;  Y : out std_logic);

end IV_24;

architecture SYN_BEHAVIORAL of IV_24 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity IV_23 is

   port( A : in std_logic;  Y : out std_logic);

end IV_23;

architecture SYN_BEHAVIORAL of IV_23 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity IV_22 is

   port( A : in std_logic;  Y : out std_logic);

end IV_22;

architecture SYN_BEHAVIORAL of IV_22 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity IV_21 is

   port( A : in std_logic;  Y : out std_logic);

end IV_21;

architecture SYN_BEHAVIORAL of IV_21 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity IV_20 is

   port( A : in std_logic;  Y : out std_logic);

end IV_20;

architecture SYN_BEHAVIORAL of IV_20 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity IV_19 is

   port( A : in std_logic;  Y : out std_logic);

end IV_19;

architecture SYN_BEHAVIORAL of IV_19 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity IV_18 is

   port( A : in std_logic;  Y : out std_logic);

end IV_18;

architecture SYN_BEHAVIORAL of IV_18 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity IV_17 is

   port( A : in std_logic;  Y : out std_logic);

end IV_17;

architecture SYN_BEHAVIORAL of IV_17 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity IV_16 is

   port( A : in std_logic;  Y : out std_logic);

end IV_16;

architecture SYN_BEHAVIORAL of IV_16 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity IV_15 is

   port( A : in std_logic;  Y : out std_logic);

end IV_15;

architecture SYN_BEHAVIORAL of IV_15 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity IV_14 is

   port( A : in std_logic;  Y : out std_logic);

end IV_14;

architecture SYN_BEHAVIORAL of IV_14 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity IV_13 is

   port( A : in std_logic;  Y : out std_logic);

end IV_13;

architecture SYN_BEHAVIORAL of IV_13 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity IV_12 is

   port( A : in std_logic;  Y : out std_logic);

end IV_12;

architecture SYN_BEHAVIORAL of IV_12 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity IV_11 is

   port( A : in std_logic;  Y : out std_logic);

end IV_11;

architecture SYN_BEHAVIORAL of IV_11 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity IV_10 is

   port( A : in std_logic;  Y : out std_logic);

end IV_10;

architecture SYN_BEHAVIORAL of IV_10 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity IV_9 is

   port( A : in std_logic;  Y : out std_logic);

end IV_9;

architecture SYN_BEHAVIORAL of IV_9 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity IV_8 is

   port( A : in std_logic;  Y : out std_logic);

end IV_8;

architecture SYN_BEHAVIORAL of IV_8 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity IV_7 is

   port( A : in std_logic;  Y : out std_logic);

end IV_7;

architecture SYN_BEHAVIORAL of IV_7 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity IV_6 is

   port( A : in std_logic;  Y : out std_logic);

end IV_6;

architecture SYN_BEHAVIORAL of IV_6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity IV_5 is

   port( A : in std_logic;  Y : out std_logic);

end IV_5;

architecture SYN_BEHAVIORAL of IV_5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity IV_4 is

   port( A : in std_logic;  Y : out std_logic);

end IV_4;

architecture SYN_BEHAVIORAL of IV_4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity IV_3 is

   port( A : in std_logic;  Y : out std_logic);

end IV_3;

architecture SYN_BEHAVIORAL of IV_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity IV_2 is

   port( A : in std_logic;  Y : out std_logic);

end IV_2;

architecture SYN_BEHAVIORAL of IV_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity IV_1 is

   port( A : in std_logic;  Y : out std_logic);

end IV_1;

architecture SYN_BEHAVIORAL of IV_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity MUX21_31 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_31;

architecture SYN_STRUCTURAL of MUX21_31 is

   component ND2_91
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_92
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_93
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_31
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_31 port map( A => S, Y => SB);
   UND1 : ND2_93 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_92 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_91 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity MUX21_30 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_30;

architecture SYN_STRUCTURAL of MUX21_30 is

   component ND2_88
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_89
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_90
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_30
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_30 port map( A => S, Y => SB);
   UND1 : ND2_90 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_89 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_88 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity MUX21_29 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_29;

architecture SYN_STRUCTURAL of MUX21_29 is

   component ND2_85
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_86
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_87
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_29
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_29 port map( A => S, Y => SB);
   UND1 : ND2_87 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_86 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_85 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity MUX21_28 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_28;

architecture SYN_STRUCTURAL of MUX21_28 is

   component ND2_82
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_83
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_84
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_28
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_28 port map( A => S, Y => SB);
   UND1 : ND2_84 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_83 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_82 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity MUX21_27 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_27;

architecture SYN_STRUCTURAL of MUX21_27 is

   component ND2_79
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_80
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_81
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_27
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_27 port map( A => S, Y => SB);
   UND1 : ND2_81 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_80 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_79 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity MUX21_26 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_26;

architecture SYN_STRUCTURAL of MUX21_26 is

   component ND2_76
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_77
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_78
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_26
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_26 port map( A => S, Y => SB);
   UND1 : ND2_78 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_77 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_76 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity MUX21_25 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_25;

architecture SYN_STRUCTURAL of MUX21_25 is

   component ND2_73
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_74
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_75
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_25
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_25 port map( A => S, Y => SB);
   UND1 : ND2_75 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_74 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_73 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity MUX21_24 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_24;

architecture SYN_STRUCTURAL of MUX21_24 is

   component ND2_70
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_71
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_72
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_24
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_24 port map( A => S, Y => SB);
   UND1 : ND2_72 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_71 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_70 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity MUX21_23 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_23;

architecture SYN_STRUCTURAL of MUX21_23 is

   component ND2_67
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_68
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_69
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_23
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_23 port map( A => S, Y => SB);
   UND1 : ND2_69 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_68 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_67 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity MUX21_22 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_22;

architecture SYN_STRUCTURAL of MUX21_22 is

   component ND2_64
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_65
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_66
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_22
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_22 port map( A => S, Y => SB);
   UND1 : ND2_66 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_65 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_64 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity MUX21_21 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_21;

architecture SYN_STRUCTURAL of MUX21_21 is

   component ND2_61
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_62
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_63
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_21
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_21 port map( A => S, Y => SB);
   UND1 : ND2_63 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_62 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_61 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity MUX21_20 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_20;

architecture SYN_STRUCTURAL of MUX21_20 is

   component ND2_58
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_59
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_60
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_20
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_20 port map( A => S, Y => SB);
   UND1 : ND2_60 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_59 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_58 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity MUX21_19 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_19;

architecture SYN_STRUCTURAL of MUX21_19 is

   component ND2_55
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_56
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_57
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_19
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_19 port map( A => S, Y => SB);
   UND1 : ND2_57 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_56 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_55 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity MUX21_18 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_18;

architecture SYN_STRUCTURAL of MUX21_18 is

   component ND2_52
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_53
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_54
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_18
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_18 port map( A => S, Y => SB);
   UND1 : ND2_54 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_53 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_52 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity MUX21_17 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_17;

architecture SYN_STRUCTURAL of MUX21_17 is

   component ND2_49
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_50
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_51
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_17
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_17 port map( A => S, Y => SB);
   UND1 : ND2_51 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_50 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_49 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity MUX21_16 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_16;

architecture SYN_STRUCTURAL of MUX21_16 is

   component ND2_46
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_47
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_48
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_16
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_16 port map( A => S, Y => SB);
   UND1 : ND2_48 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_47 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_46 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity MUX21_15 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_15;

architecture SYN_STRUCTURAL of MUX21_15 is

   component ND2_43
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_44
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_45
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_15
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_15 port map( A => S, Y => SB);
   UND1 : ND2_45 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_44 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_43 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity MUX21_14 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_14;

architecture SYN_STRUCTURAL of MUX21_14 is

   component ND2_40
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_41
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_42
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_14
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_14 port map( A => S, Y => SB);
   UND1 : ND2_42 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_41 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_40 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity MUX21_13 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_13;

architecture SYN_STRUCTURAL of MUX21_13 is

   component ND2_37
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_38
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_39
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_13
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_13 port map( A => S, Y => SB);
   UND1 : ND2_39 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_38 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_37 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity MUX21_12 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_12;

architecture SYN_STRUCTURAL of MUX21_12 is

   component ND2_34
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_35
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_36
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_12
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_12 port map( A => S, Y => SB);
   UND1 : ND2_36 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_35 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_34 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity MUX21_11 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_11;

architecture SYN_STRUCTURAL of MUX21_11 is

   component ND2_31
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_32
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_33
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_11
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_11 port map( A => S, Y => SB);
   UND1 : ND2_33 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_32 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_31 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity MUX21_10 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_10;

architecture SYN_STRUCTURAL of MUX21_10 is

   component ND2_28
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_29
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_30
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_10
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_10 port map( A => S, Y => SB);
   UND1 : ND2_30 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_29 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_28 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity MUX21_9 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_9;

architecture SYN_STRUCTURAL of MUX21_9 is

   component ND2_25
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_26
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_27
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_9
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_9 port map( A => S, Y => SB);
   UND1 : ND2_27 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_26 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_25 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity MUX21_8 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_8;

architecture SYN_STRUCTURAL of MUX21_8 is

   component ND2_22
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_23
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_24
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_8
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_8 port map( A => S, Y => SB);
   UND1 : ND2_24 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_23 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_22 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity MUX21_7 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_7;

architecture SYN_STRUCTURAL of MUX21_7 is

   component ND2_19
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_20
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_21
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_7
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_7 port map( A => S, Y => SB);
   UND1 : ND2_21 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_20 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_19 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity MUX21_6 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_6;

architecture SYN_STRUCTURAL of MUX21_6 is

   component ND2_16
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_17
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_18
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_6
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_6 port map( A => S, Y => SB);
   UND1 : ND2_18 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_17 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_16 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity MUX21_5 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_5;

architecture SYN_STRUCTURAL of MUX21_5 is

   component ND2_13
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_14
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_15
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_5
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_5 port map( A => S, Y => SB);
   UND1 : ND2_15 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_14 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_13 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity MUX21_4 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_4;

architecture SYN_STRUCTURAL of MUX21_4 is

   component ND2_10
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_11
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_12
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_4 port map( A => S, Y => SB);
   UND1 : ND2_12 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_11 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_10 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity MUX21_3 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_3;

architecture SYN_STRUCTURAL of MUX21_3 is

   component ND2_7
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_8
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_9
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_3
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_3 port map( A => S, Y => SB);
   UND1 : ND2_9 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_8 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_7 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity MUX21_2 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_2;

architecture SYN_STRUCTURAL of MUX21_2 is

   component ND2_4
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_5
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_6
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_2 port map( A => S, Y => SB);
   UND1 : ND2_6 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_5 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_4 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity MUX21_1 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_1;

architecture SYN_STRUCTURAL of MUX21_1 is

   component ND2_1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_3
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_1 port map( A => S, Y => SB);
   UND1 : ND2_3 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_2 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_1 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity FA_63 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_63;

architecture SYN_Behavioural of FA_63 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => c_in, B => n11, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => c_out);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n11, B2 => c_in, ZN => n10);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity FA_62 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_62;

architecture SYN_Behavioural of FA_62 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => c_in, B => n11, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => c_out);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n11, B2 => c_in, ZN => n10);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity FA_61 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_61;

architecture SYN_Behavioural of FA_61 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => c_in, B => n11, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => c_out);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n11, B2 => c_in, ZN => n10);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity FA_60 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_60;

architecture SYN_Behavioural of FA_60 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => c_in, B => n11, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => c_out);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n11, B2 => c_in, ZN => n10);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity FA_59 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_59;

architecture SYN_Behavioural of FA_59 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => c_in, B => n11, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => c_out);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n11, B2 => c_in, ZN => n10);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity FA_58 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_58;

architecture SYN_Behavioural of FA_58 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => c_in, B => n11, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => c_out);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n11, B2 => c_in, ZN => n10);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity FA_57 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_57;

architecture SYN_Behavioural of FA_57 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => c_in, B => n11, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => c_out);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n11, B2 => c_in, ZN => n10);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity FA_56 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_56;

architecture SYN_Behavioural of FA_56 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => c_in, B => n11, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => c_out);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n11, B2 => c_in, ZN => n10);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity FA_55 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_55;

architecture SYN_Behavioural of FA_55 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => c_in, B => n11, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => c_out);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n11, B2 => c_in, ZN => n10);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity FA_54 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_54;

architecture SYN_Behavioural of FA_54 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => c_in, B => n11, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => c_out);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n11, B2 => c_in, ZN => n10);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity FA_53 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_53;

architecture SYN_Behavioural of FA_53 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => c_in, B => n11, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => c_out);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n11, B2 => c_in, ZN => n10);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity FA_52 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_52;

architecture SYN_Behavioural of FA_52 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => c_in, B => n11, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => c_out);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n11, B2 => c_in, ZN => n10);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity FA_51 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_51;

architecture SYN_Behavioural of FA_51 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => c_in, B => n11, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => c_out);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n11, B2 => c_in, ZN => n10);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity FA_50 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_50;

architecture SYN_Behavioural of FA_50 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => c_in, B => n11, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => c_out);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n11, B2 => c_in, ZN => n10);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity FA_49 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_49;

architecture SYN_Behavioural of FA_49 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => c_in, B => n11, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => c_out);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n11, B2 => c_in, ZN => n10);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity FA_48 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_48;

architecture SYN_Behavioural of FA_48 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => c_in, B => n11, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => c_out);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n11, B2 => c_in, ZN => n10);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity FA_47 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_47;

architecture SYN_Behavioural of FA_47 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => c_in, B => n11, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => c_out);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n11, B2 => c_in, ZN => n10);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity FA_46 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_46;

architecture SYN_Behavioural of FA_46 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => c_in, B => n11, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => c_out);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n11, B2 => c_in, ZN => n10);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity FA_45 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_45;

architecture SYN_Behavioural of FA_45 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => c_in, B => n11, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => c_out);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n11, B2 => c_in, ZN => n10);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity FA_44 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_44;

architecture SYN_Behavioural of FA_44 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => c_in, B => n11, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => c_out);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n11, B2 => c_in, ZN => n10);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity FA_43 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_43;

architecture SYN_Behavioural of FA_43 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => c_in, B => n11, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => c_out);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n11, B2 => c_in, ZN => n10);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity FA_42 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_42;

architecture SYN_Behavioural of FA_42 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => c_in, B => n11, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => c_out);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n11, B2 => c_in, ZN => n10);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity FA_41 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_41;

architecture SYN_Behavioural of FA_41 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => c_in, B => n11, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => c_out);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n11, B2 => c_in, ZN => n10);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity FA_40 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_40;

architecture SYN_Behavioural of FA_40 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => c_in, B => n11, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => c_out);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n11, B2 => c_in, ZN => n10);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity FA_39 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_39;

architecture SYN_Behavioural of FA_39 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => c_in, B => n11, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => c_out);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n11, B2 => c_in, ZN => n10);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity FA_38 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_38;

architecture SYN_Behavioural of FA_38 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => c_in, B => n11, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => c_out);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n11, B2 => c_in, ZN => n10);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity FA_37 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_37;

architecture SYN_Behavioural of FA_37 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => c_in, B => n11, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => c_out);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n11, B2 => c_in, ZN => n10);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity FA_36 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_36;

architecture SYN_Behavioural of FA_36 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => c_in, B => n11, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => c_out);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n11, B2 => c_in, ZN => n10);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity FA_35 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_35;

architecture SYN_Behavioural of FA_35 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => c_in, B => n11, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => c_out);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n11, B2 => c_in, ZN => n10);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity FA_34 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_34;

architecture SYN_Behavioural of FA_34 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => c_in, B => n11, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => c_out);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n11, B2 => c_in, ZN => n10);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity FA_33 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_33;

architecture SYN_Behavioural of FA_33 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => c_in, B => n11, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => c_out);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n11, B2 => c_in, ZN => n10);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity FA_32 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_32;

architecture SYN_Behavioural of FA_32 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => c_in, B => n11, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => c_out);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n11, B2 => c_in, ZN => n10);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity FA_31 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_31;

architecture SYN_Behavioural of FA_31 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => c_in, B => n11, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => c_out);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n11, B2 => c_in, ZN => n10);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity FA_30 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_30;

architecture SYN_Behavioural of FA_30 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => c_in, B => n11, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => c_out);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n11, B2 => c_in, ZN => n10);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity FA_29 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_29;

architecture SYN_Behavioural of FA_29 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => c_in, B => n11, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => c_out);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n11, B2 => c_in, ZN => n10);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity FA_28 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_28;

architecture SYN_Behavioural of FA_28 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => c_in, B => n11, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => c_out);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n11, B2 => c_in, ZN => n10);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity FA_27 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_27;

architecture SYN_Behavioural of FA_27 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => c_in, B => n11, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => c_out);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n11, B2 => c_in, ZN => n10);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity FA_26 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_26;

architecture SYN_Behavioural of FA_26 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => c_in, B => n11, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => c_out);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n11, B2 => c_in, ZN => n10);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity FA_25 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_25;

architecture SYN_Behavioural of FA_25 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => c_in, B => n11, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => c_out);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n11, B2 => c_in, ZN => n10);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity FA_24 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_24;

architecture SYN_Behavioural of FA_24 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => c_in, B => n11, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => c_out);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n11, B2 => c_in, ZN => n10);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity FA_23 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_23;

architecture SYN_Behavioural of FA_23 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => c_in, B => n11, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => c_out);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n11, B2 => c_in, ZN => n10);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity FA_22 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_22;

architecture SYN_Behavioural of FA_22 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => c_in, B => n11, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => c_out);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n11, B2 => c_in, ZN => n10);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity FA_21 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_21;

architecture SYN_Behavioural of FA_21 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => c_in, B => n11, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => c_out);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n11, B2 => c_in, ZN => n10);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity FA_20 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_20;

architecture SYN_Behavioural of FA_20 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => c_in, B => n11, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => c_out);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n11, B2 => c_in, ZN => n10);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity FA_19 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_19;

architecture SYN_Behavioural of FA_19 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => c_in, B => n11, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => c_out);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n11, B2 => c_in, ZN => n10);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity FA_18 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_18;

architecture SYN_Behavioural of FA_18 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => c_in, B => n11, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => c_out);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n11, B2 => c_in, ZN => n10);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity FA_17 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_17;

architecture SYN_Behavioural of FA_17 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => c_in, B => n11, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => c_out);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n11, B2 => c_in, ZN => n10);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity FA_16 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_16;

architecture SYN_Behavioural of FA_16 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => c_in, B => n11, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => c_out);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n11, B2 => c_in, ZN => n10);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity FA_15 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_15;

architecture SYN_Behavioural of FA_15 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => c_in, B => n11, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => c_out);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n11, B2 => c_in, ZN => n10);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity FA_14 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_14;

architecture SYN_Behavioural of FA_14 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => c_in, B => n11, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => c_out);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n11, B2 => c_in, ZN => n10);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity FA_13 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_13;

architecture SYN_Behavioural of FA_13 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => c_in, B => n11, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => c_out);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n11, B2 => c_in, ZN => n10);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity FA_12 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_12;

architecture SYN_Behavioural of FA_12 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => c_in, B => n11, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => c_out);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n11, B2 => c_in, ZN => n10);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity FA_11 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_11;

architecture SYN_Behavioural of FA_11 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => c_in, B => n11, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => c_out);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n11, B2 => c_in, ZN => n10);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity FA_10 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_10;

architecture SYN_Behavioural of FA_10 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => c_in, B => n11, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => c_out);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n11, B2 => c_in, ZN => n10);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity FA_9 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_9;

architecture SYN_Behavioural of FA_9 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => c_in, B => n11, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => c_out);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n11, B2 => c_in, ZN => n10);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity FA_8 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_8;

architecture SYN_Behavioural of FA_8 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => c_in, B => n11, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => c_out);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n11, B2 => c_in, ZN => n10);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity FA_7 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_7;

architecture SYN_Behavioural of FA_7 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => c_in, B => n11, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => c_out);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n11, B2 => c_in, ZN => n10);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity FA_6 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_6;

architecture SYN_Behavioural of FA_6 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => c_in, B => n11, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => c_out);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n11, B2 => c_in, ZN => n10);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity FA_5 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_5;

architecture SYN_Behavioural of FA_5 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => c_in, B => n11, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => c_out);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n11, B2 => c_in, ZN => n10);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity FA_4 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_4;

architecture SYN_Behavioural of FA_4 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => c_in, B => n11, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => c_out);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n11, B2 => c_in, ZN => n10);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity FA_3 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_3;

architecture SYN_Behavioural of FA_3 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => c_in, B => n11, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => c_out);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n11, B2 => c_in, ZN => n10);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity FA_2 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_2;

architecture SYN_Behavioural of FA_2 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => c_in, B => n11, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => c_out);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n11, B2 => c_in, ZN => n10);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity FA_1 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_1;

architecture SYN_Behavioural of FA_1 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => c_in, B => n11, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => c_out);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n11, B2 => c_in, ZN => n10);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity MUX21_GENERIC_NBIT4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_7;

architecture SYN_STRUCTURAL of MUX21_GENERIC_NBIT4_7 is

   component MUX21_25
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_26
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_27
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_28
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUX21GENI_0 : MUX21_28 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUX21GENI_1 : MUX21_27 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUX21GENI_2 : MUX21_26 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUX21GENI_3 : MUX21_25 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity MUX21_GENERIC_NBIT4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_6;

architecture SYN_STRUCTURAL of MUX21_GENERIC_NBIT4_6 is

   component MUX21_21
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_22
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_23
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_24
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUX21GENI_0 : MUX21_24 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUX21GENI_1 : MUX21_23 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUX21GENI_2 : MUX21_22 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUX21GENI_3 : MUX21_21 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity MUX21_GENERIC_NBIT4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_5;

architecture SYN_STRUCTURAL of MUX21_GENERIC_NBIT4_5 is

   component MUX21_17
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_18
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_19
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_20
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUX21GENI_0 : MUX21_20 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUX21GENI_1 : MUX21_19 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUX21GENI_2 : MUX21_18 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUX21GENI_3 : MUX21_17 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity MUX21_GENERIC_NBIT4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_4;

architecture SYN_STRUCTURAL of MUX21_GENERIC_NBIT4_4 is

   component MUX21_13
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_14
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_15
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_16
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUX21GENI_0 : MUX21_16 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUX21GENI_1 : MUX21_15 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUX21GENI_2 : MUX21_14 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUX21GENI_3 : MUX21_13 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity MUX21_GENERIC_NBIT4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_3;

architecture SYN_STRUCTURAL of MUX21_GENERIC_NBIT4_3 is

   component MUX21_9
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_10
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_11
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_12
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUX21GENI_0 : MUX21_12 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUX21GENI_1 : MUX21_11 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUX21GENI_2 : MUX21_10 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUX21GENI_3 : MUX21_9 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity MUX21_GENERIC_NBIT4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_2;

architecture SYN_STRUCTURAL of MUX21_GENERIC_NBIT4_2 is

   component MUX21_5
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_6
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_7
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_8
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUX21GENI_0 : MUX21_8 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUX21GENI_1 : MUX21_7 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUX21GENI_2 : MUX21_6 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUX21GENI_3 : MUX21_5 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity MUX21_GENERIC_NBIT4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_1;

architecture SYN_STRUCTURAL of MUX21_GENERIC_NBIT4_1 is

   component MUX21_1
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_2
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_3
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_4
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUX21GENI_0 : MUX21_4 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUX21GENI_1 : MUX21_3 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUX21GENI_2 : MUX21_2 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUX21GENI_3 : MUX21_1 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity RCA_size4_15 is

   port( a, b : in std_logic_vector (3 downto 0);  c_in : in std_logic;  c_out 
         : out std_logic;  sum : out std_logic_vector (3 downto 0));

end RCA_size4_15;

architecture SYN_Structural of RCA_size4_15 is

   component FA_57
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_58
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_59
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_60
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   signal temp_3_port, temp_2_port, temp_1_port : std_logic;

begin
   
   fa_i_0 : FA_60 port map( a => a(0), b => b(0), c_in => c_in, c_out => 
                           temp_1_port, s => sum(0));
   fa_i_1 : FA_59 port map( a => a(1), b => b(1), c_in => temp_1_port, c_out =>
                           temp_2_port, s => sum(1));
   fa_i_2 : FA_58 port map( a => a(2), b => b(2), c_in => temp_2_port, c_out =>
                           temp_3_port, s => sum(2));
   fa_i_3 : FA_57 port map( a => a(3), b => b(3), c_in => temp_3_port, c_out =>
                           c_out, s => sum(3));

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity RCA_size4_14 is

   port( a, b : in std_logic_vector (3 downto 0);  c_in : in std_logic;  c_out 
         : out std_logic;  sum : out std_logic_vector (3 downto 0));

end RCA_size4_14;

architecture SYN_Structural of RCA_size4_14 is

   component FA_53
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_54
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_55
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_56
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   signal temp_3_port, temp_2_port, temp_1_port : std_logic;

begin
   
   fa_i_0 : FA_56 port map( a => a(0), b => b(0), c_in => c_in, c_out => 
                           temp_1_port, s => sum(0));
   fa_i_1 : FA_55 port map( a => a(1), b => b(1), c_in => temp_1_port, c_out =>
                           temp_2_port, s => sum(1));
   fa_i_2 : FA_54 port map( a => a(2), b => b(2), c_in => temp_2_port, c_out =>
                           temp_3_port, s => sum(2));
   fa_i_3 : FA_53 port map( a => a(3), b => b(3), c_in => temp_3_port, c_out =>
                           c_out, s => sum(3));

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity RCA_size4_13 is

   port( a, b : in std_logic_vector (3 downto 0);  c_in : in std_logic;  c_out 
         : out std_logic;  sum : out std_logic_vector (3 downto 0));

end RCA_size4_13;

architecture SYN_Structural of RCA_size4_13 is

   component FA_49
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_50
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_51
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_52
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   signal temp_3_port, temp_2_port, temp_1_port : std_logic;

begin
   
   fa_i_0 : FA_52 port map( a => a(0), b => b(0), c_in => c_in, c_out => 
                           temp_1_port, s => sum(0));
   fa_i_1 : FA_51 port map( a => a(1), b => b(1), c_in => temp_1_port, c_out =>
                           temp_2_port, s => sum(1));
   fa_i_2 : FA_50 port map( a => a(2), b => b(2), c_in => temp_2_port, c_out =>
                           temp_3_port, s => sum(2));
   fa_i_3 : FA_49 port map( a => a(3), b => b(3), c_in => temp_3_port, c_out =>
                           c_out, s => sum(3));

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity RCA_size4_12 is

   port( a, b : in std_logic_vector (3 downto 0);  c_in : in std_logic;  c_out 
         : out std_logic;  sum : out std_logic_vector (3 downto 0));

end RCA_size4_12;

architecture SYN_Structural of RCA_size4_12 is

   component FA_45
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_46
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_47
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_48
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   signal temp_3_port, temp_2_port, temp_1_port : std_logic;

begin
   
   fa_i_0 : FA_48 port map( a => a(0), b => b(0), c_in => c_in, c_out => 
                           temp_1_port, s => sum(0));
   fa_i_1 : FA_47 port map( a => a(1), b => b(1), c_in => temp_1_port, c_out =>
                           temp_2_port, s => sum(1));
   fa_i_2 : FA_46 port map( a => a(2), b => b(2), c_in => temp_2_port, c_out =>
                           temp_3_port, s => sum(2));
   fa_i_3 : FA_45 port map( a => a(3), b => b(3), c_in => temp_3_port, c_out =>
                           c_out, s => sum(3));

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity RCA_size4_11 is

   port( a, b : in std_logic_vector (3 downto 0);  c_in : in std_logic;  c_out 
         : out std_logic;  sum : out std_logic_vector (3 downto 0));

end RCA_size4_11;

architecture SYN_Structural of RCA_size4_11 is

   component FA_41
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_42
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_43
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_44
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   signal temp_3_port, temp_2_port, temp_1_port : std_logic;

begin
   
   fa_i_0 : FA_44 port map( a => a(0), b => b(0), c_in => c_in, c_out => 
                           temp_1_port, s => sum(0));
   fa_i_1 : FA_43 port map( a => a(1), b => b(1), c_in => temp_1_port, c_out =>
                           temp_2_port, s => sum(1));
   fa_i_2 : FA_42 port map( a => a(2), b => b(2), c_in => temp_2_port, c_out =>
                           temp_3_port, s => sum(2));
   fa_i_3 : FA_41 port map( a => a(3), b => b(3), c_in => temp_3_port, c_out =>
                           c_out, s => sum(3));

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity RCA_size4_10 is

   port( a, b : in std_logic_vector (3 downto 0);  c_in : in std_logic;  c_out 
         : out std_logic;  sum : out std_logic_vector (3 downto 0));

end RCA_size4_10;

architecture SYN_Structural of RCA_size4_10 is

   component FA_37
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_38
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_39
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_40
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   signal temp_3_port, temp_2_port, temp_1_port : std_logic;

begin
   
   fa_i_0 : FA_40 port map( a => a(0), b => b(0), c_in => c_in, c_out => 
                           temp_1_port, s => sum(0));
   fa_i_1 : FA_39 port map( a => a(1), b => b(1), c_in => temp_1_port, c_out =>
                           temp_2_port, s => sum(1));
   fa_i_2 : FA_38 port map( a => a(2), b => b(2), c_in => temp_2_port, c_out =>
                           temp_3_port, s => sum(2));
   fa_i_3 : FA_37 port map( a => a(3), b => b(3), c_in => temp_3_port, c_out =>
                           c_out, s => sum(3));

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity RCA_size4_9 is

   port( a, b : in std_logic_vector (3 downto 0);  c_in : in std_logic;  c_out 
         : out std_logic;  sum : out std_logic_vector (3 downto 0));

end RCA_size4_9;

architecture SYN_Structural of RCA_size4_9 is

   component FA_33
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_34
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_35
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_36
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   signal temp_3_port, temp_2_port, temp_1_port : std_logic;

begin
   
   fa_i_0 : FA_36 port map( a => a(0), b => b(0), c_in => c_in, c_out => 
                           temp_1_port, s => sum(0));
   fa_i_1 : FA_35 port map( a => a(1), b => b(1), c_in => temp_1_port, c_out =>
                           temp_2_port, s => sum(1));
   fa_i_2 : FA_34 port map( a => a(2), b => b(2), c_in => temp_2_port, c_out =>
                           temp_3_port, s => sum(2));
   fa_i_3 : FA_33 port map( a => a(3), b => b(3), c_in => temp_3_port, c_out =>
                           c_out, s => sum(3));

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity RCA_size4_8 is

   port( a, b : in std_logic_vector (3 downto 0);  c_in : in std_logic;  c_out 
         : out std_logic;  sum : out std_logic_vector (3 downto 0));

end RCA_size4_8;

architecture SYN_Structural of RCA_size4_8 is

   component FA_29
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_30
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_31
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_32
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   signal temp_3_port, temp_2_port, temp_1_port : std_logic;

begin
   
   fa_i_0 : FA_32 port map( a => a(0), b => b(0), c_in => c_in, c_out => 
                           temp_1_port, s => sum(0));
   fa_i_1 : FA_31 port map( a => a(1), b => b(1), c_in => temp_1_port, c_out =>
                           temp_2_port, s => sum(1));
   fa_i_2 : FA_30 port map( a => a(2), b => b(2), c_in => temp_2_port, c_out =>
                           temp_3_port, s => sum(2));
   fa_i_3 : FA_29 port map( a => a(3), b => b(3), c_in => temp_3_port, c_out =>
                           c_out, s => sum(3));

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity RCA_size4_7 is

   port( a, b : in std_logic_vector (3 downto 0);  c_in : in std_logic;  c_out 
         : out std_logic;  sum : out std_logic_vector (3 downto 0));

end RCA_size4_7;

architecture SYN_Structural of RCA_size4_7 is

   component FA_25
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_26
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_27
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_28
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   signal temp_3_port, temp_2_port, temp_1_port : std_logic;

begin
   
   fa_i_0 : FA_28 port map( a => a(0), b => b(0), c_in => c_in, c_out => 
                           temp_1_port, s => sum(0));
   fa_i_1 : FA_27 port map( a => a(1), b => b(1), c_in => temp_1_port, c_out =>
                           temp_2_port, s => sum(1));
   fa_i_2 : FA_26 port map( a => a(2), b => b(2), c_in => temp_2_port, c_out =>
                           temp_3_port, s => sum(2));
   fa_i_3 : FA_25 port map( a => a(3), b => b(3), c_in => temp_3_port, c_out =>
                           c_out, s => sum(3));

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity RCA_size4_6 is

   port( a, b : in std_logic_vector (3 downto 0);  c_in : in std_logic;  c_out 
         : out std_logic;  sum : out std_logic_vector (3 downto 0));

end RCA_size4_6;

architecture SYN_Structural of RCA_size4_6 is

   component FA_21
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_22
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_23
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_24
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   signal temp_3_port, temp_2_port, temp_1_port : std_logic;

begin
   
   fa_i_0 : FA_24 port map( a => a(0), b => b(0), c_in => c_in, c_out => 
                           temp_1_port, s => sum(0));
   fa_i_1 : FA_23 port map( a => a(1), b => b(1), c_in => temp_1_port, c_out =>
                           temp_2_port, s => sum(1));
   fa_i_2 : FA_22 port map( a => a(2), b => b(2), c_in => temp_2_port, c_out =>
                           temp_3_port, s => sum(2));
   fa_i_3 : FA_21 port map( a => a(3), b => b(3), c_in => temp_3_port, c_out =>
                           c_out, s => sum(3));

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity RCA_size4_5 is

   port( a, b : in std_logic_vector (3 downto 0);  c_in : in std_logic;  c_out 
         : out std_logic;  sum : out std_logic_vector (3 downto 0));

end RCA_size4_5;

architecture SYN_Structural of RCA_size4_5 is

   component FA_17
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_18
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_19
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_20
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   signal temp_3_port, temp_2_port, temp_1_port : std_logic;

begin
   
   fa_i_0 : FA_20 port map( a => a(0), b => b(0), c_in => c_in, c_out => 
                           temp_1_port, s => sum(0));
   fa_i_1 : FA_19 port map( a => a(1), b => b(1), c_in => temp_1_port, c_out =>
                           temp_2_port, s => sum(1));
   fa_i_2 : FA_18 port map( a => a(2), b => b(2), c_in => temp_2_port, c_out =>
                           temp_3_port, s => sum(2));
   fa_i_3 : FA_17 port map( a => a(3), b => b(3), c_in => temp_3_port, c_out =>
                           c_out, s => sum(3));

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity RCA_size4_4 is

   port( a, b : in std_logic_vector (3 downto 0);  c_in : in std_logic;  c_out 
         : out std_logic;  sum : out std_logic_vector (3 downto 0));

end RCA_size4_4;

architecture SYN_Structural of RCA_size4_4 is

   component FA_13
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_14
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_15
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_16
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   signal temp_3_port, temp_2_port, temp_1_port : std_logic;

begin
   
   fa_i_0 : FA_16 port map( a => a(0), b => b(0), c_in => c_in, c_out => 
                           temp_1_port, s => sum(0));
   fa_i_1 : FA_15 port map( a => a(1), b => b(1), c_in => temp_1_port, c_out =>
                           temp_2_port, s => sum(1));
   fa_i_2 : FA_14 port map( a => a(2), b => b(2), c_in => temp_2_port, c_out =>
                           temp_3_port, s => sum(2));
   fa_i_3 : FA_13 port map( a => a(3), b => b(3), c_in => temp_3_port, c_out =>
                           c_out, s => sum(3));

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity RCA_size4_3 is

   port( a, b : in std_logic_vector (3 downto 0);  c_in : in std_logic;  c_out 
         : out std_logic;  sum : out std_logic_vector (3 downto 0));

end RCA_size4_3;

architecture SYN_Structural of RCA_size4_3 is

   component FA_9
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_10
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_11
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_12
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   signal temp_3_port, temp_2_port, temp_1_port : std_logic;

begin
   
   fa_i_0 : FA_12 port map( a => a(0), b => b(0), c_in => c_in, c_out => 
                           temp_1_port, s => sum(0));
   fa_i_1 : FA_11 port map( a => a(1), b => b(1), c_in => temp_1_port, c_out =>
                           temp_2_port, s => sum(1));
   fa_i_2 : FA_10 port map( a => a(2), b => b(2), c_in => temp_2_port, c_out =>
                           temp_3_port, s => sum(2));
   fa_i_3 : FA_9 port map( a => a(3), b => b(3), c_in => temp_3_port, c_out => 
                           c_out, s => sum(3));

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity RCA_size4_2 is

   port( a, b : in std_logic_vector (3 downto 0);  c_in : in std_logic;  c_out 
         : out std_logic;  sum : out std_logic_vector (3 downto 0));

end RCA_size4_2;

architecture SYN_Structural of RCA_size4_2 is

   component FA_5
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_6
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_7
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_8
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   signal temp_3_port, temp_2_port, temp_1_port : std_logic;

begin
   
   fa_i_0 : FA_8 port map( a => a(0), b => b(0), c_in => c_in, c_out => 
                           temp_1_port, s => sum(0));
   fa_i_1 : FA_7 port map( a => a(1), b => b(1), c_in => temp_1_port, c_out => 
                           temp_2_port, s => sum(1));
   fa_i_2 : FA_6 port map( a => a(2), b => b(2), c_in => temp_2_port, c_out => 
                           temp_3_port, s => sum(2));
   fa_i_3 : FA_5 port map( a => a(3), b => b(3), c_in => temp_3_port, c_out => 
                           c_out, s => sum(3));

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity RCA_size4_1 is

   port( a, b : in std_logic_vector (3 downto 0);  c_in : in std_logic;  c_out 
         : out std_logic;  sum : out std_logic_vector (3 downto 0));

end RCA_size4_1;

architecture SYN_Structural of RCA_size4_1 is

   component FA_1
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_2
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_3
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_4
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   signal temp_3_port, temp_2_port, temp_1_port : std_logic;

begin
   
   fa_i_0 : FA_4 port map( a => a(0), b => b(0), c_in => c_in, c_out => 
                           temp_1_port, s => sum(0));
   fa_i_1 : FA_3 port map( a => a(1), b => b(1), c_in => temp_1_port, c_out => 
                           temp_2_port, s => sum(1));
   fa_i_2 : FA_2 port map( a => a(2), b => b(2), c_in => temp_2_port, c_out => 
                           temp_3_port, s => sum(2));
   fa_i_3 : FA_1 port map( a => a(3), b => b(3), c_in => temp_3_port, c_out => 
                           c_out, s => sum(3));

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity SUM_BLOCK_K4_7 is

   port( a, b : in std_logic_vector (3 downto 0);  C_gen : in std_logic;  sum :
         out std_logic_vector (3 downto 0));

end SUM_BLOCK_K4_7;

architecture SYN_Structural of SUM_BLOCK_K4_7 is

   component MUX21_GENERIC_NBIT4_7
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_size4_13
      port( a, b : in std_logic_vector (3 downto 0);  c_in : in std_logic;  
            c_out : out std_logic;  sum : out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_size4_14
      port( a, b : in std_logic_vector (3 downto 0);  c_in : in std_logic;  
            c_out : out std_logic;  sum : out std_logic_vector (3 downto 0));
   end component;
   
   signal X_Logic1_port, X_Logic0_port, SUM1_3_port, SUM1_2_port, SUM1_1_port, 
      SUM1_0_port, SUM2_3_port, SUM2_2_port, SUM2_1_port, SUM2_0_port, n_1000, 
      n_1001 : std_logic;

begin
   
   RCA_CIN0 : RCA_size4_14 port map( a(3) => a(3), a(2) => a(2), a(1) => a(1), 
                           a(0) => a(0), b(3) => b(3), b(2) => b(2), b(1) => 
                           b(1), b(0) => b(0), c_in => X_Logic0_port, c_out => 
                           n_1000, sum(3) => SUM1_3_port, sum(2) => SUM1_2_port
                           , sum(1) => SUM1_1_port, sum(0) => SUM1_0_port);
   RCA_CIN1 : RCA_size4_13 port map( a(3) => a(3), a(2) => a(2), a(1) => a(1), 
                           a(0) => a(0), b(3) => b(3), b(2) => b(2), b(1) => 
                           b(1), b(0) => b(0), c_in => X_Logic1_port, c_out => 
                           n_1001, sum(3) => SUM2_3_port, sum(2) => SUM2_2_port
                           , sum(1) => SUM2_1_port, sum(0) => SUM2_0_port);
   MPX : MUX21_GENERIC_NBIT4_7 port map( A(3) => SUM2_3_port, A(2) => 
                           SUM2_2_port, A(1) => SUM2_1_port, A(0) => 
                           SUM2_0_port, B(3) => SUM1_3_port, B(2) => 
                           SUM1_2_port, B(1) => SUM1_1_port, B(0) => 
                           SUM1_0_port, SEL => C_gen, Y(3) => sum(3), Y(2) => 
                           sum(2), Y(1) => sum(1), Y(0) => sum(0));
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity SUM_BLOCK_K4_6 is

   port( a, b : in std_logic_vector (3 downto 0);  C_gen : in std_logic;  sum :
         out std_logic_vector (3 downto 0));

end SUM_BLOCK_K4_6;

architecture SYN_Structural of SUM_BLOCK_K4_6 is

   component MUX21_GENERIC_NBIT4_6
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_size4_11
      port( a, b : in std_logic_vector (3 downto 0);  c_in : in std_logic;  
            c_out : out std_logic;  sum : out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_size4_12
      port( a, b : in std_logic_vector (3 downto 0);  c_in : in std_logic;  
            c_out : out std_logic;  sum : out std_logic_vector (3 downto 0));
   end component;
   
   signal X_Logic1_port, X_Logic0_port, SUM1_3_port, SUM1_2_port, SUM1_1_port, 
      SUM1_0_port, SUM2_3_port, SUM2_2_port, SUM2_1_port, SUM2_0_port, n_1002, 
      n_1003 : std_logic;

begin
   
   RCA_CIN0 : RCA_size4_12 port map( a(3) => a(3), a(2) => a(2), a(1) => a(1), 
                           a(0) => a(0), b(3) => b(3), b(2) => b(2), b(1) => 
                           b(1), b(0) => b(0), c_in => X_Logic0_port, c_out => 
                           n_1002, sum(3) => SUM1_3_port, sum(2) => SUM1_2_port
                           , sum(1) => SUM1_1_port, sum(0) => SUM1_0_port);
   RCA_CIN1 : RCA_size4_11 port map( a(3) => a(3), a(2) => a(2), a(1) => a(1), 
                           a(0) => a(0), b(3) => b(3), b(2) => b(2), b(1) => 
                           b(1), b(0) => b(0), c_in => X_Logic1_port, c_out => 
                           n_1003, sum(3) => SUM2_3_port, sum(2) => SUM2_2_port
                           , sum(1) => SUM2_1_port, sum(0) => SUM2_0_port);
   MPX : MUX21_GENERIC_NBIT4_6 port map( A(3) => SUM2_3_port, A(2) => 
                           SUM2_2_port, A(1) => SUM2_1_port, A(0) => 
                           SUM2_0_port, B(3) => SUM1_3_port, B(2) => 
                           SUM1_2_port, B(1) => SUM1_1_port, B(0) => 
                           SUM1_0_port, SEL => C_gen, Y(3) => sum(3), Y(2) => 
                           sum(2), Y(1) => sum(1), Y(0) => sum(0));
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity SUM_BLOCK_K4_5 is

   port( a, b : in std_logic_vector (3 downto 0);  C_gen : in std_logic;  sum :
         out std_logic_vector (3 downto 0));

end SUM_BLOCK_K4_5;

architecture SYN_Structural of SUM_BLOCK_K4_5 is

   component MUX21_GENERIC_NBIT4_5
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_size4_9
      port( a, b : in std_logic_vector (3 downto 0);  c_in : in std_logic;  
            c_out : out std_logic;  sum : out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_size4_10
      port( a, b : in std_logic_vector (3 downto 0);  c_in : in std_logic;  
            c_out : out std_logic;  sum : out std_logic_vector (3 downto 0));
   end component;
   
   signal X_Logic1_port, X_Logic0_port, SUM1_3_port, SUM1_2_port, SUM1_1_port, 
      SUM1_0_port, SUM2_3_port, SUM2_2_port, SUM2_1_port, SUM2_0_port, n_1004, 
      n_1005 : std_logic;

begin
   
   RCA_CIN0 : RCA_size4_10 port map( a(3) => a(3), a(2) => a(2), a(1) => a(1), 
                           a(0) => a(0), b(3) => b(3), b(2) => b(2), b(1) => 
                           b(1), b(0) => b(0), c_in => X_Logic0_port, c_out => 
                           n_1004, sum(3) => SUM1_3_port, sum(2) => SUM1_2_port
                           , sum(1) => SUM1_1_port, sum(0) => SUM1_0_port);
   RCA_CIN1 : RCA_size4_9 port map( a(3) => a(3), a(2) => a(2), a(1) => a(1), 
                           a(0) => a(0), b(3) => b(3), b(2) => b(2), b(1) => 
                           b(1), b(0) => b(0), c_in => X_Logic1_port, c_out => 
                           n_1005, sum(3) => SUM2_3_port, sum(2) => SUM2_2_port
                           , sum(1) => SUM2_1_port, sum(0) => SUM2_0_port);
   MPX : MUX21_GENERIC_NBIT4_5 port map( A(3) => SUM2_3_port, A(2) => 
                           SUM2_2_port, A(1) => SUM2_1_port, A(0) => 
                           SUM2_0_port, B(3) => SUM1_3_port, B(2) => 
                           SUM1_2_port, B(1) => SUM1_1_port, B(0) => 
                           SUM1_0_port, SEL => C_gen, Y(3) => sum(3), Y(2) => 
                           sum(2), Y(1) => sum(1), Y(0) => sum(0));
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity SUM_BLOCK_K4_4 is

   port( a, b : in std_logic_vector (3 downto 0);  C_gen : in std_logic;  sum :
         out std_logic_vector (3 downto 0));

end SUM_BLOCK_K4_4;

architecture SYN_Structural of SUM_BLOCK_K4_4 is

   component MUX21_GENERIC_NBIT4_4
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_size4_7
      port( a, b : in std_logic_vector (3 downto 0);  c_in : in std_logic;  
            c_out : out std_logic;  sum : out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_size4_8
      port( a, b : in std_logic_vector (3 downto 0);  c_in : in std_logic;  
            c_out : out std_logic;  sum : out std_logic_vector (3 downto 0));
   end component;
   
   signal X_Logic1_port, X_Logic0_port, SUM1_3_port, SUM1_2_port, SUM1_1_port, 
      SUM1_0_port, SUM2_3_port, SUM2_2_port, SUM2_1_port, SUM2_0_port, n_1006, 
      n_1007 : std_logic;

begin
   
   RCA_CIN0 : RCA_size4_8 port map( a(3) => a(3), a(2) => a(2), a(1) => a(1), 
                           a(0) => a(0), b(3) => b(3), b(2) => b(2), b(1) => 
                           b(1), b(0) => b(0), c_in => X_Logic0_port, c_out => 
                           n_1006, sum(3) => SUM1_3_port, sum(2) => SUM1_2_port
                           , sum(1) => SUM1_1_port, sum(0) => SUM1_0_port);
   RCA_CIN1 : RCA_size4_7 port map( a(3) => a(3), a(2) => a(2), a(1) => a(1), 
                           a(0) => a(0), b(3) => b(3), b(2) => b(2), b(1) => 
                           b(1), b(0) => b(0), c_in => X_Logic1_port, c_out => 
                           n_1007, sum(3) => SUM2_3_port, sum(2) => SUM2_2_port
                           , sum(1) => SUM2_1_port, sum(0) => SUM2_0_port);
   MPX : MUX21_GENERIC_NBIT4_4 port map( A(3) => SUM2_3_port, A(2) => 
                           SUM2_2_port, A(1) => SUM2_1_port, A(0) => 
                           SUM2_0_port, B(3) => SUM1_3_port, B(2) => 
                           SUM1_2_port, B(1) => SUM1_1_port, B(0) => 
                           SUM1_0_port, SEL => C_gen, Y(3) => sum(3), Y(2) => 
                           sum(2), Y(1) => sum(1), Y(0) => sum(0));
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity SUM_BLOCK_K4_3 is

   port( a, b : in std_logic_vector (3 downto 0);  C_gen : in std_logic;  sum :
         out std_logic_vector (3 downto 0));

end SUM_BLOCK_K4_3;

architecture SYN_Structural of SUM_BLOCK_K4_3 is

   component MUX21_GENERIC_NBIT4_3
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_size4_5
      port( a, b : in std_logic_vector (3 downto 0);  c_in : in std_logic;  
            c_out : out std_logic;  sum : out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_size4_6
      port( a, b : in std_logic_vector (3 downto 0);  c_in : in std_logic;  
            c_out : out std_logic;  sum : out std_logic_vector (3 downto 0));
   end component;
   
   signal X_Logic1_port, X_Logic0_port, SUM1_3_port, SUM1_2_port, SUM1_1_port, 
      SUM1_0_port, SUM2_3_port, SUM2_2_port, SUM2_1_port, SUM2_0_port, n_1008, 
      n_1009 : std_logic;

begin
   
   RCA_CIN0 : RCA_size4_6 port map( a(3) => a(3), a(2) => a(2), a(1) => a(1), 
                           a(0) => a(0), b(3) => b(3), b(2) => b(2), b(1) => 
                           b(1), b(0) => b(0), c_in => X_Logic0_port, c_out => 
                           n_1008, sum(3) => SUM1_3_port, sum(2) => SUM1_2_port
                           , sum(1) => SUM1_1_port, sum(0) => SUM1_0_port);
   RCA_CIN1 : RCA_size4_5 port map( a(3) => a(3), a(2) => a(2), a(1) => a(1), 
                           a(0) => a(0), b(3) => b(3), b(2) => b(2), b(1) => 
                           b(1), b(0) => b(0), c_in => X_Logic1_port, c_out => 
                           n_1009, sum(3) => SUM2_3_port, sum(2) => SUM2_2_port
                           , sum(1) => SUM2_1_port, sum(0) => SUM2_0_port);
   MPX : MUX21_GENERIC_NBIT4_3 port map( A(3) => SUM2_3_port, A(2) => 
                           SUM2_2_port, A(1) => SUM2_1_port, A(0) => 
                           SUM2_0_port, B(3) => SUM1_3_port, B(2) => 
                           SUM1_2_port, B(1) => SUM1_1_port, B(0) => 
                           SUM1_0_port, SEL => C_gen, Y(3) => sum(3), Y(2) => 
                           sum(2), Y(1) => sum(1), Y(0) => sum(0));
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity SUM_BLOCK_K4_2 is

   port( a, b : in std_logic_vector (3 downto 0);  C_gen : in std_logic;  sum :
         out std_logic_vector (3 downto 0));

end SUM_BLOCK_K4_2;

architecture SYN_Structural of SUM_BLOCK_K4_2 is

   component MUX21_GENERIC_NBIT4_2
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_size4_3
      port( a, b : in std_logic_vector (3 downto 0);  c_in : in std_logic;  
            c_out : out std_logic;  sum : out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_size4_4
      port( a, b : in std_logic_vector (3 downto 0);  c_in : in std_logic;  
            c_out : out std_logic;  sum : out std_logic_vector (3 downto 0));
   end component;
   
   signal X_Logic1_port, X_Logic0_port, SUM1_3_port, SUM1_2_port, SUM1_1_port, 
      SUM1_0_port, SUM2_3_port, SUM2_2_port, SUM2_1_port, SUM2_0_port, n_1010, 
      n_1011 : std_logic;

begin
   
   RCA_CIN0 : RCA_size4_4 port map( a(3) => a(3), a(2) => a(2), a(1) => a(1), 
                           a(0) => a(0), b(3) => b(3), b(2) => b(2), b(1) => 
                           b(1), b(0) => b(0), c_in => X_Logic0_port, c_out => 
                           n_1010, sum(3) => SUM1_3_port, sum(2) => SUM1_2_port
                           , sum(1) => SUM1_1_port, sum(0) => SUM1_0_port);
   RCA_CIN1 : RCA_size4_3 port map( a(3) => a(3), a(2) => a(2), a(1) => a(1), 
                           a(0) => a(0), b(3) => b(3), b(2) => b(2), b(1) => 
                           b(1), b(0) => b(0), c_in => X_Logic1_port, c_out => 
                           n_1011, sum(3) => SUM2_3_port, sum(2) => SUM2_2_port
                           , sum(1) => SUM2_1_port, sum(0) => SUM2_0_port);
   MPX : MUX21_GENERIC_NBIT4_2 port map( A(3) => SUM2_3_port, A(2) => 
                           SUM2_2_port, A(1) => SUM2_1_port, A(0) => 
                           SUM2_0_port, B(3) => SUM1_3_port, B(2) => 
                           SUM1_2_port, B(1) => SUM1_1_port, B(0) => 
                           SUM1_0_port, SEL => C_gen, Y(3) => sum(3), Y(2) => 
                           sum(2), Y(1) => sum(1), Y(0) => sum(0));
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity SUM_BLOCK_K4_1 is

   port( a, b : in std_logic_vector (3 downto 0);  C_gen : in std_logic;  sum :
         out std_logic_vector (3 downto 0));

end SUM_BLOCK_K4_1;

architecture SYN_Structural of SUM_BLOCK_K4_1 is

   component MUX21_GENERIC_NBIT4_1
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_size4_1
      port( a, b : in std_logic_vector (3 downto 0);  c_in : in std_logic;  
            c_out : out std_logic;  sum : out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_size4_2
      port( a, b : in std_logic_vector (3 downto 0);  c_in : in std_logic;  
            c_out : out std_logic;  sum : out std_logic_vector (3 downto 0));
   end component;
   
   signal X_Logic1_port, X_Logic0_port, SUM1_3_port, SUM1_2_port, SUM1_1_port, 
      SUM1_0_port, SUM2_3_port, SUM2_2_port, SUM2_1_port, SUM2_0_port, n_1012, 
      n_1013 : std_logic;

begin
   
   RCA_CIN0 : RCA_size4_2 port map( a(3) => a(3), a(2) => a(2), a(1) => a(1), 
                           a(0) => a(0), b(3) => b(3), b(2) => b(2), b(1) => 
                           b(1), b(0) => b(0), c_in => X_Logic0_port, c_out => 
                           n_1012, sum(3) => SUM1_3_port, sum(2) => SUM1_2_port
                           , sum(1) => SUM1_1_port, sum(0) => SUM1_0_port);
   RCA_CIN1 : RCA_size4_1 port map( a(3) => a(3), a(2) => a(2), a(1) => a(1), 
                           a(0) => a(0), b(3) => b(3), b(2) => b(2), b(1) => 
                           b(1), b(0) => b(0), c_in => X_Logic1_port, c_out => 
                           n_1013, sum(3) => SUM2_3_port, sum(2) => SUM2_2_port
                           , sum(1) => SUM2_1_port, sum(0) => SUM2_0_port);
   MPX : MUX21_GENERIC_NBIT4_1 port map( A(3) => SUM2_3_port, A(2) => 
                           SUM2_2_port, A(1) => SUM2_1_port, A(0) => 
                           SUM2_0_port, B(3) => SUM1_3_port, B(2) => 
                           SUM1_2_port, B(1) => SUM1_1_port, B(0) => 
                           SUM1_0_port, SEL => C_gen, Y(3) => sum(3), Y(2) => 
                           sum(2), Y(1) => sum(1), Y(0) => sum(0));
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity PG_BLOCK_26 is

   port( PIK, GIK, PK1J, GK1J : in std_logic;  GIJ, PIJ : out std_logic);

end PG_BLOCK_26;

architecture SYN_Behavioral of PG_BLOCK_26 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PK1J, A2 => PIK, ZN => PIJ);
   U2 : INV_X1 port map( A => n7, ZN => GIJ);
   U3 : AOI21_X1 port map( B1 => PIK, B2 => GK1J, A => GIK, ZN => n7);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity PG_BLOCK_25 is

   port( PIK, GIK, PK1J, GK1J : in std_logic;  GIJ, PIJ : out std_logic);

end PG_BLOCK_25;

architecture SYN_Behavioral of PG_BLOCK_25 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => PIK, Z => n7);
   U2 : INV_X1 port map( A => n8, ZN => GIJ);
   U3 : AOI21_X1 port map( B1 => PIK, B2 => GK1J, A => GIK, ZN => n8);
   U4 : AND2_X1 port map( A1 => n7, A2 => PK1J, ZN => PIJ);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity PG_BLOCK_24 is

   port( PIK, GIK, PK1J, GK1J : in std_logic;  GIJ, PIJ : out std_logic);

end PG_BLOCK_24;

architecture SYN_Behavioral of PG_BLOCK_24 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => PIK, B2 => GK1J, A => GIK, ZN => n7);
   U2 : AND2_X1 port map( A1 => PK1J, A2 => PIK, ZN => PIJ);
   U3 : INV_X1 port map( A => n7, ZN => GIJ);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity PG_BLOCK_23 is

   port( PIK, GIK, PK1J, GK1J : in std_logic;  GIJ, PIJ : out std_logic);

end PG_BLOCK_23;

architecture SYN_Behavioral of PG_BLOCK_23 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PK1J, A2 => PIK, ZN => PIJ);
   U2 : INV_X1 port map( A => n7, ZN => GIJ);
   U3 : AOI21_X1 port map( B1 => PIK, B2 => GK1J, A => GIK, ZN => n7);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity PG_BLOCK_22 is

   port( PIK, GIK, PK1J, GK1J : in std_logic;  GIJ, PIJ : out std_logic);

end PG_BLOCK_22;

architecture SYN_Behavioral of PG_BLOCK_22 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PK1J, A2 => PIK, ZN => PIJ);
   U2 : INV_X1 port map( A => n7, ZN => GIJ);
   U3 : AOI21_X1 port map( B1 => PIK, B2 => GK1J, A => GIK, ZN => n7);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity PG_BLOCK_21 is

   port( PIK, GIK, PK1J, GK1J : in std_logic;  GIJ, PIJ : out std_logic);

end PG_BLOCK_21;

architecture SYN_Behavioral of PG_BLOCK_21 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n7, ZN => GIJ);
   U2 : AND2_X1 port map( A1 => PIK, A2 => PK1J, ZN => PIJ);
   U3 : AOI21_X1 port map( B1 => PIK, B2 => GK1J, A => GIK, ZN => n7);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity PG_BLOCK_20 is

   port( PIK, GIK, PK1J, GK1J : in std_logic;  GIJ, PIJ : out std_logic);

end PG_BLOCK_20;

architecture SYN_Behavioral of PG_BLOCK_20 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n7, ZN => GIJ);
   U2 : AOI21_X1 port map( B1 => PIK, B2 => GK1J, A => GIK, ZN => n7);
   U3 : AND2_X1 port map( A1 => PK1J, A2 => PIK, ZN => PIJ);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity PG_BLOCK_19 is

   port( PIK, GIK, PK1J, GK1J : in std_logic;  GIJ, PIJ : out std_logic);

end PG_BLOCK_19;

architecture SYN_Behavioral of PG_BLOCK_19 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PK1J, A2 => PIK, ZN => PIJ);
   U2 : INV_X1 port map( A => n7, ZN => GIJ);
   U3 : AOI21_X1 port map( B1 => PIK, B2 => GK1J, A => GIK, ZN => n7);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity PG_BLOCK_18 is

   port( PIK, GIK, PK1J, GK1J : in std_logic;  GIJ, PIJ : out std_logic);

end PG_BLOCK_18;

architecture SYN_Behavioral of PG_BLOCK_18 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n7, ZN => GIJ);
   U2 : AOI21_X1 port map( B1 => PIK, B2 => GK1J, A => GIK, ZN => n7);
   U3 : AND2_X1 port map( A1 => PK1J, A2 => PIK, ZN => PIJ);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity PG_BLOCK_17 is

   port( PIK, GIK, PK1J, GK1J : in std_logic;  GIJ, PIJ : out std_logic);

end PG_BLOCK_17;

architecture SYN_Behavioral of PG_BLOCK_17 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n7, ZN => GIJ);
   U2 : AOI21_X1 port map( B1 => PIK, B2 => GK1J, A => GIK, ZN => n7);
   U3 : AND2_X1 port map( A1 => PIK, A2 => PK1J, ZN => PIJ);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity PG_BLOCK_16 is

   port( PIK, GIK, PK1J, GK1J : in std_logic;  GIJ, PIJ : out std_logic);

end PG_BLOCK_16;

architecture SYN_Behavioral of PG_BLOCK_16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n7, ZN => GIJ);
   U2 : AOI21_X1 port map( B1 => PIK, B2 => GK1J, A => GIK, ZN => n7);
   U3 : AND2_X1 port map( A1 => PK1J, A2 => PIK, ZN => PIJ);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity PG_BLOCK_15 is

   port( PIK, GIK, PK1J, GK1J : in std_logic;  GIJ, PIJ : out std_logic);

end PG_BLOCK_15;

architecture SYN_Behavioral of PG_BLOCK_15 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n7, ZN => GIJ);
   U2 : AOI21_X1 port map( B1 => PIK, B2 => GK1J, A => GIK, ZN => n7);
   U3 : AND2_X1 port map( A1 => PK1J, A2 => PIK, ZN => PIJ);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity PG_BLOCK_14 is

   port( PIK, GIK, PK1J, GK1J : in std_logic;  GIJ, PIJ : out std_logic);

end PG_BLOCK_14;

architecture SYN_Behavioral of PG_BLOCK_14 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n7, ZN => GIJ);
   U2 : AOI21_X1 port map( B1 => PIK, B2 => GK1J, A => GIK, ZN => n7);
   U3 : AND2_X1 port map( A1 => PK1J, A2 => PIK, ZN => PIJ);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity PG_BLOCK_13 is

   port( PIK, GIK, PK1J, GK1J : in std_logic;  GIJ, PIJ : out std_logic);

end PG_BLOCK_13;

architecture SYN_Behavioral of PG_BLOCK_13 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n7, ZN => GIJ);
   U2 : AOI21_X1 port map( B1 => PIK, B2 => GK1J, A => GIK, ZN => n7);
   U3 : AND2_X1 port map( A1 => PK1J, A2 => PIK, ZN => PIJ);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity PG_BLOCK_12 is

   port( PIK, GIK, PK1J, GK1J : in std_logic;  GIJ, PIJ : out std_logic);

end PG_BLOCK_12;

architecture SYN_Behavioral of PG_BLOCK_12 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PK1J, A2 => PIK, ZN => PIJ);
   U2 : INV_X1 port map( A => n7, ZN => GIJ);
   U3 : AOI21_X1 port map( B1 => PIK, B2 => GK1J, A => GIK, ZN => n7);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity PG_BLOCK_11 is

   port( PIK, GIK, PK1J, GK1J : in std_logic;  GIJ, PIJ : out std_logic);

end PG_BLOCK_11;

architecture SYN_Behavioral of PG_BLOCK_11 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PK1J, A2 => PIK, ZN => PIJ);
   U2 : AOI21_X1 port map( B1 => PIK, B2 => GK1J, A => GIK, ZN => n7);
   U3 : INV_X1 port map( A => n7, ZN => GIJ);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity PG_BLOCK_10 is

   port( PIK, GIK, PK1J, GK1J : in std_logic;  GIJ, PIJ : out std_logic);

end PG_BLOCK_10;

architecture SYN_Behavioral of PG_BLOCK_10 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PK1J, A2 => PIK, ZN => PIJ);
   U2 : AOI21_X1 port map( B1 => PIK, B2 => GK1J, A => GIK, ZN => n7);
   U3 : INV_X1 port map( A => n7, ZN => GIJ);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity PG_BLOCK_9 is

   port( PIK, GIK, PK1J, GK1J : in std_logic;  GIJ, PIJ : out std_logic);

end PG_BLOCK_9;

architecture SYN_Behavioral of PG_BLOCK_9 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => PIK, B2 => GK1J, A => GIK, ZN => n7);
   U2 : AND2_X1 port map( A1 => PK1J, A2 => PIK, ZN => PIJ);
   U3 : INV_X1 port map( A => n7, ZN => GIJ);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity PG_BLOCK_8 is

   port( PIK, GIK, PK1J, GK1J : in std_logic;  GIJ, PIJ : out std_logic);

end PG_BLOCK_8;

architecture SYN_Behavioral of PG_BLOCK_8 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => PIK, B2 => GK1J, A => GIK, ZN => n7);
   U2 : AND2_X1 port map( A1 => PK1J, A2 => PIK, ZN => PIJ);
   U3 : INV_X1 port map( A => n7, ZN => GIJ);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity PG_BLOCK_7 is

   port( PIK, GIK, PK1J, GK1J : in std_logic;  GIJ, PIJ : out std_logic);

end PG_BLOCK_7;

architecture SYN_Behavioral of PG_BLOCK_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n7, ZN => GIJ);
   U2 : AOI21_X1 port map( B1 => PIK, B2 => GK1J, A => GIK, ZN => n7);
   U3 : AND2_X1 port map( A1 => PK1J, A2 => PIK, ZN => PIJ);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity PG_BLOCK_6 is

   port( PIK, GIK, PK1J, GK1J : in std_logic;  GIJ, PIJ : out std_logic);

end PG_BLOCK_6;

architecture SYN_Behavioral of PG_BLOCK_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n7, ZN => GIJ);
   U2 : AOI21_X1 port map( B1 => PIK, B2 => GK1J, A => GIK, ZN => n7);
   U3 : AND2_X1 port map( A1 => PK1J, A2 => PIK, ZN => PIJ);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity PG_BLOCK_5 is

   port( PIK, GIK, PK1J, GK1J : in std_logic;  GIJ, PIJ : out std_logic);

end PG_BLOCK_5;

architecture SYN_Behavioral of PG_BLOCK_5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PK1J, A2 => PIK, ZN => PIJ);
   U2 : AOI21_X1 port map( B1 => GK1J, B2 => PIK, A => GIK, ZN => n7);
   U3 : INV_X1 port map( A => n7, ZN => GIJ);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity PG_BLOCK_4 is

   port( PIK, GIK, PK1J, GK1J : in std_logic;  GIJ, PIJ : out std_logic);

end PG_BLOCK_4;

architecture SYN_Behavioral of PG_BLOCK_4 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PK1J, A2 => PIK, ZN => PIJ);
   U2 : INV_X1 port map( A => n7, ZN => GIJ);
   U3 : AOI21_X1 port map( B1 => PIK, B2 => GK1J, A => GIK, ZN => n7);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity PG_BLOCK_3 is

   port( PIK, GIK, PK1J, GK1J : in std_logic;  GIJ, PIJ : out std_logic);

end PG_BLOCK_3;

architecture SYN_Behavioral of PG_BLOCK_3 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n7, ZN => GIJ);
   U2 : AOI21_X1 port map( B1 => PIK, B2 => GK1J, A => GIK, ZN => n7);
   U3 : AND2_X1 port map( A1 => PK1J, A2 => PIK, ZN => PIJ);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity PG_BLOCK_2 is

   port( PIK, GIK, PK1J, GK1J : in std_logic;  GIJ, PIJ : out std_logic);

end PG_BLOCK_2;

architecture SYN_Behavioral of PG_BLOCK_2 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PK1J, A2 => PIK, ZN => PIJ);
   U2 : INV_X1 port map( A => n7, ZN => GIJ);
   U3 : AOI21_X1 port map( B1 => GK1J, B2 => PIK, A => GIK, ZN => n7);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity PG_BLOCK_1 is

   port( PIK, GIK, PK1J, GK1J : in std_logic;  GIJ, PIJ : out std_logic);

end PG_BLOCK_1;

architecture SYN_Behavioral of PG_BLOCK_1 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PK1J, A2 => PIK, ZN => PIJ);
   U2 : INV_X1 port map( A => n7, ZN => GIJ);
   U3 : AOI21_X1 port map( B1 => PIK, B2 => GK1J, A => GIK, ZN => n7);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity G_BLOCK_8 is

   port( PIK, GIK, GK1J : in std_logic;  GIJ : out std_logic);

end G_BLOCK_8;

architecture SYN_Behavioral of G_BLOCK_8 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => PIK, B2 => GK1J, A => GIK, ZN => n7);
   U2 : INV_X1 port map( A => n7, ZN => GIJ);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity G_BLOCK_7 is

   port( PIK, GIK, GK1J : in std_logic;  GIJ : out std_logic);

end G_BLOCK_7;

architecture SYN_Behavioral of G_BLOCK_7 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n7, ZN => GIJ);
   U2 : AOI21_X1 port map( B1 => PIK, B2 => GK1J, A => GIK, ZN => n7);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity G_BLOCK_6 is

   port( PIK, GIK, GK1J : in std_logic;  GIJ : out std_logic);

end G_BLOCK_6;

architecture SYN_Behavioral of G_BLOCK_6 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n7, ZN => GIJ);
   U2 : AOI21_X1 port map( B1 => PIK, B2 => GK1J, A => GIK, ZN => n7);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity G_BLOCK_5 is

   port( PIK, GIK, GK1J : in std_logic;  GIJ : out std_logic);

end G_BLOCK_5;

architecture SYN_Behavioral of G_BLOCK_5 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => GIK, ZN => n7);
   U2 : NAND2_X1 port map( A1 => n7, A2 => n8, ZN => GIJ);
   U3 : NAND2_X1 port map( A1 => GK1J, A2 => PIK, ZN => n8);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity G_BLOCK_4 is

   port( PIK, GIK, GK1J : in std_logic;  GIJ : out std_logic);

end G_BLOCK_4;

architecture SYN_Behavioral of G_BLOCK_4 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => GIK, ZN => n7);
   U2 : NAND2_X2 port map( A1 => n7, A2 => n8, ZN => GIJ);
   U3 : NAND2_X1 port map( A1 => GK1J, A2 => PIK, ZN => n8);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity G_BLOCK_3 is

   port( PIK, GIK, GK1J : in std_logic;  GIJ : out std_logic);

end G_BLOCK_3;

architecture SYN_Behavioral of G_BLOCK_3 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => GIK, ZN => n7);
   U2 : NAND2_X2 port map( A1 => n7, A2 => n8, ZN => GIJ);
   U3 : NAND2_X1 port map( A1 => GK1J, A2 => PIK, ZN => n8);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity G_BLOCK_2 is

   port( PIK, GIK, GK1J : in std_logic;  GIJ : out std_logic);

end G_BLOCK_2;

architecture SYN_Behavioral of G_BLOCK_2 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => GIK, ZN => n7);
   U2 : NAND2_X2 port map( A1 => n7, A2 => n8, ZN => GIJ);
   U3 : NAND2_X1 port map( A1 => GK1J, A2 => PIK, ZN => n8);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity G_BLOCK_1 is

   port( PIK, GIK, GK1J : in std_logic;  GIJ : out std_logic);

end G_BLOCK_1;

architecture SYN_Behavioral of G_BLOCK_1 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n7, ZN => GIJ);
   U2 : AOI21_X1 port map( B1 => PIK, B2 => GK1J, A => GIK, ZN => n7);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity PG_NET_31 is

   port( A, B : in std_logic;  P, G : out std_logic);

end PG_NET_31;

architecture SYN_Behavioral of PG_NET_31 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity PG_NET_30 is

   port( A, B : in std_logic;  P, G : out std_logic);

end PG_NET_30;

architecture SYN_Behavioral of PG_NET_30 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity PG_NET_29 is

   port( A, B : in std_logic;  P, G : out std_logic);

end PG_NET_29;

architecture SYN_Behavioral of PG_NET_29 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity PG_NET_28 is

   port( A, B : in std_logic;  P, G : out std_logic);

end PG_NET_28;

architecture SYN_Behavioral of PG_NET_28 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity PG_NET_27 is

   port( A, B : in std_logic;  P, G : out std_logic);

end PG_NET_27;

architecture SYN_Behavioral of PG_NET_27 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity PG_NET_26 is

   port( A, B : in std_logic;  P, G : out std_logic);

end PG_NET_26;

architecture SYN_Behavioral of PG_NET_26 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity PG_NET_25 is

   port( A, B : in std_logic;  P, G : out std_logic);

end PG_NET_25;

architecture SYN_Behavioral of PG_NET_25 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity PG_NET_24 is

   port( A, B : in std_logic;  P, G : out std_logic);

end PG_NET_24;

architecture SYN_Behavioral of PG_NET_24 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity PG_NET_23 is

   port( A, B : in std_logic;  P, G : out std_logic);

end PG_NET_23;

architecture SYN_Behavioral of PG_NET_23 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity PG_NET_22 is

   port( A, B : in std_logic;  P, G : out std_logic);

end PG_NET_22;

architecture SYN_Behavioral of PG_NET_22 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity PG_NET_21 is

   port( A, B : in std_logic;  P, G : out std_logic);

end PG_NET_21;

architecture SYN_Behavioral of PG_NET_21 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => n2, ZN => n3);
   U2 : NAND2_X1 port map( A1 => n1, A2 => A, ZN => n4);
   U3 : NAND2_X1 port map( A1 => n3, A2 => n4, ZN => P);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : INV_X1 port map( A => A, ZN => n2);
   U6 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity PG_NET_20 is

   port( A, B : in std_logic;  P, G : out std_logic);

end PG_NET_20;

architecture SYN_Behavioral of PG_NET_20 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity PG_NET_19 is

   port( A, B : in std_logic;  P, G : out std_logic);

end PG_NET_19;

architecture SYN_Behavioral of PG_NET_19 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity PG_NET_18 is

   port( A, B : in std_logic;  P, G : out std_logic);

end PG_NET_18;

architecture SYN_Behavioral of PG_NET_18 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity PG_NET_17 is

   port( A, B : in std_logic;  P, G : out std_logic);

end PG_NET_17;

architecture SYN_Behavioral of PG_NET_17 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n2, A2 => B, ZN => n3);
   U2 : NAND2_X1 port map( A1 => n1, A2 => A, ZN => n4);
   U3 : NAND2_X1 port map( A1 => n3, A2 => n4, ZN => P);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : INV_X1 port map( A => A, ZN => n2);
   U6 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity PG_NET_16 is

   port( A, B : in std_logic;  P, G : out std_logic);

end PG_NET_16;

architecture SYN_Behavioral of PG_NET_16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity PG_NET_15 is

   port( A, B : in std_logic;  P, G : out std_logic);

end PG_NET_15;

architecture SYN_Behavioral of PG_NET_15 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity PG_NET_14 is

   port( A, B : in std_logic;  P, G : out std_logic);

end PG_NET_14;

architecture SYN_Behavioral of PG_NET_14 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity PG_NET_13 is

   port( A, B : in std_logic;  P, G : out std_logic);

end PG_NET_13;

architecture SYN_Behavioral of PG_NET_13 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity PG_NET_12 is

   port( A, B : in std_logic;  P, G : out std_logic);

end PG_NET_12;

architecture SYN_Behavioral of PG_NET_12 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity PG_NET_11 is

   port( A, B : in std_logic;  P, G : out std_logic);

end PG_NET_11;

architecture SYN_Behavioral of PG_NET_11 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity PG_NET_10 is

   port( A, B : in std_logic;  P, G : out std_logic);

end PG_NET_10;

architecture SYN_Behavioral of PG_NET_10 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity PG_NET_9 is

   port( A, B : in std_logic;  P, G : out std_logic);

end PG_NET_9;

architecture SYN_Behavioral of PG_NET_9 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n2, A2 => B, ZN => n3);
   U2 : NAND2_X1 port map( A1 => n1, A2 => A, ZN => n4);
   U3 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => P);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : INV_X1 port map( A => A, ZN => n2);
   U6 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity PG_NET_8 is

   port( A, B : in std_logic;  P, G : out std_logic);

end PG_NET_8;

architecture SYN_Behavioral of PG_NET_8 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity PG_NET_7 is

   port( A, B : in std_logic;  P, G : out std_logic);

end PG_NET_7;

architecture SYN_Behavioral of PG_NET_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity PG_NET_6 is

   port( A, B : in std_logic;  P, G : out std_logic);

end PG_NET_6;

architecture SYN_Behavioral of PG_NET_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity PG_NET_5 is

   port( A, B : in std_logic;  P, G : out std_logic);

end PG_NET_5;

architecture SYN_Behavioral of PG_NET_5 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity PG_NET_4 is

   port( A, B : in std_logic;  P, G : out std_logic);

end PG_NET_4;

architecture SYN_Behavioral of PG_NET_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity PG_NET_3 is

   port( A, B : in std_logic;  P, G : out std_logic);

end PG_NET_3;

architecture SYN_Behavioral of PG_NET_3 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity PG_NET_2 is

   port( A, B : in std_logic;  P, G : out std_logic);

end PG_NET_2;

architecture SYN_Behavioral of PG_NET_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity PG_NET_1 is

   port( A, B : in std_logic;  P, G : out std_logic);

end PG_NET_1;

architecture SYN_Behavioral of PG_NET_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity ND2_0 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_0;

architecture SYN_ARCH2 of ND2_0 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity IV_0 is

   port( A : in std_logic;  Y : out std_logic);

end IV_0;

architecture SYN_BEHAVIORAL of IV_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity MUX21_0 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_0;

architecture SYN_STRUCTURAL of MUX21_0 is

   component ND2_94
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_95
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_0
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_0
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_0 port map( A => S, Y => SB);
   UND1 : ND2_0 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_95 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_94 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity FA_0 is

   port( a, b, c_in : in std_logic;  c_out, s : out std_logic);

end FA_0;

architecture SYN_Behavioural of FA_0 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => c_in, B => n2, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => c_out);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n2, B2 => c_in, ZN => n3);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity MUX21_GENERIC_NBIT4_0 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_0;

architecture SYN_STRUCTURAL of MUX21_GENERIC_NBIT4_0 is

   component MUX21_29
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_30
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_31
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_0
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUX21GENI_0 : MUX21_0 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUX21GENI_1 : MUX21_31 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUX21GENI_2 : MUX21_30 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUX21GENI_3 : MUX21_29 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity RCA_size4_0 is

   port( a, b : in std_logic_vector (3 downto 0);  c_in : in std_logic;  c_out 
         : out std_logic;  sum : out std_logic_vector (3 downto 0));

end RCA_size4_0;

architecture SYN_Structural of RCA_size4_0 is

   component FA_61
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_62
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_63
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   component FA_0
      port( a, b, c_in : in std_logic;  c_out, s : out std_logic);
   end component;
   
   signal temp_3_port, temp_2_port, temp_1_port : std_logic;

begin
   
   fa_i_0 : FA_0 port map( a => a(0), b => b(0), c_in => c_in, c_out => 
                           temp_1_port, s => sum(0));
   fa_i_1 : FA_63 port map( a => a(1), b => b(1), c_in => temp_1_port, c_out =>
                           temp_2_port, s => sum(1));
   fa_i_2 : FA_62 port map( a => a(2), b => b(2), c_in => temp_2_port, c_out =>
                           temp_3_port, s => sum(2));
   fa_i_3 : FA_61 port map( a => a(3), b => b(3), c_in => temp_3_port, c_out =>
                           c_out, s => sum(3));

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity SUM_BLOCK_K4_0 is

   port( a, b : in std_logic_vector (3 downto 0);  C_gen : in std_logic;  sum :
         out std_logic_vector (3 downto 0));

end SUM_BLOCK_K4_0;

architecture SYN_Structural of SUM_BLOCK_K4_0 is

   component MUX21_GENERIC_NBIT4_0
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_size4_15
      port( a, b : in std_logic_vector (3 downto 0);  c_in : in std_logic;  
            c_out : out std_logic;  sum : out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_size4_0
      port( a, b : in std_logic_vector (3 downto 0);  c_in : in std_logic;  
            c_out : out std_logic;  sum : out std_logic_vector (3 downto 0));
   end component;
   
   signal X_Logic1_port, X_Logic0_port, SUM1_3_port, SUM1_2_port, SUM1_1_port, 
      SUM1_0_port, SUM2_3_port, SUM2_2_port, SUM2_1_port, SUM2_0_port, n_1014, 
      n_1015 : std_logic;

begin
   
   RCA_CIN0 : RCA_size4_0 port map( a(3) => a(3), a(2) => a(2), a(1) => a(1), 
                           a(0) => a(0), b(3) => b(3), b(2) => b(2), b(1) => 
                           b(1), b(0) => b(0), c_in => X_Logic0_port, c_out => 
                           n_1014, sum(3) => SUM1_3_port, sum(2) => SUM1_2_port
                           , sum(1) => SUM1_1_port, sum(0) => SUM1_0_port);
   RCA_CIN1 : RCA_size4_15 port map( a(3) => a(3), a(2) => a(2), a(1) => a(1), 
                           a(0) => a(0), b(3) => b(3), b(2) => b(2), b(1) => 
                           b(1), b(0) => b(0), c_in => X_Logic1_port, c_out => 
                           n_1015, sum(3) => SUM2_3_port, sum(2) => SUM2_2_port
                           , sum(1) => SUM2_1_port, sum(0) => SUM2_0_port);
   MPX : MUX21_GENERIC_NBIT4_0 port map( A(3) => SUM2_3_port, A(2) => 
                           SUM2_2_port, A(1) => SUM2_1_port, A(0) => 
                           SUM2_0_port, B(3) => SUM1_3_port, B(2) => 
                           SUM1_2_port, B(1) => SUM1_1_port, B(0) => 
                           SUM1_0_port, SEL => C_gen, Y(3) => sum(3), Y(2) => 
                           sum(2), Y(1) => sum(1), Y(0) => sum(0));
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity PG_BLOCK_0 is

   port( PIK, GIK, PK1J, GK1J : in std_logic;  GIJ, PIJ : out std_logic);

end PG_BLOCK_0;

architecture SYN_Behavioral of PG_BLOCK_0 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => GIJ);
   U2 : AND2_X1 port map( A1 => PK1J, A2 => PIK, ZN => PIJ);
   U3 : AOI21_X1 port map( B1 => PIK, B2 => GK1J, A => GIK, ZN => n2);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity G_BLOCK_0 is

   port( PIK, GIK, GK1J : in std_logic;  GIJ : out std_logic);

end G_BLOCK_0;

architecture SYN_Behavioral of G_BLOCK_0 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => GIJ);
   U2 : AOI21_X1 port map( B1 => PIK, B2 => GK1J, A => GIK, ZN => n2);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity PG_NET_0 is

   port( A, B : in std_logic;  P, G : out std_logic);

end PG_NET_0;

architecture SYN_Behavioral of PG_NET_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity SUM_GENERATOR_N32_K4 is

   port( carries : in std_logic_vector (7 downto 0);  A, B : in 
         std_logic_vector (31 downto 0);  SUM : out std_logic_vector (31 downto
         0));

end SUM_GENERATOR_N32_K4;

architecture SYN_Structural of SUM_GENERATOR_N32_K4 is

   component SUM_BLOCK_K4_1
      port( a, b : in std_logic_vector (3 downto 0);  C_gen : in std_logic;  
            sum : out std_logic_vector (3 downto 0));
   end component;
   
   component SUM_BLOCK_K4_2
      port( a, b : in std_logic_vector (3 downto 0);  C_gen : in std_logic;  
            sum : out std_logic_vector (3 downto 0));
   end component;
   
   component SUM_BLOCK_K4_3
      port( a, b : in std_logic_vector (3 downto 0);  C_gen : in std_logic;  
            sum : out std_logic_vector (3 downto 0));
   end component;
   
   component SUM_BLOCK_K4_4
      port( a, b : in std_logic_vector (3 downto 0);  C_gen : in std_logic;  
            sum : out std_logic_vector (3 downto 0));
   end component;
   
   component SUM_BLOCK_K4_5
      port( a, b : in std_logic_vector (3 downto 0);  C_gen : in std_logic;  
            sum : out std_logic_vector (3 downto 0));
   end component;
   
   component SUM_BLOCK_K4_6
      port( a, b : in std_logic_vector (3 downto 0);  C_gen : in std_logic;  
            sum : out std_logic_vector (3 downto 0));
   end component;
   
   component SUM_BLOCK_K4_7
      port( a, b : in std_logic_vector (3 downto 0);  C_gen : in std_logic;  
            sum : out std_logic_vector (3 downto 0));
   end component;
   
   component SUM_BLOCK_K4_0
      port( a, b : in std_logic_vector (3 downto 0);  C_gen : in std_logic;  
            sum : out std_logic_vector (3 downto 0));
   end component;

begin
   
   SBi_0 : SUM_BLOCK_K4_0 port map( a(3) => A(3), a(2) => A(2), a(1) => A(1), 
                           a(0) => A(0), b(3) => B(3), b(2) => B(2), b(1) => 
                           B(1), b(0) => B(0), C_gen => carries(0), sum(3) => 
                           SUM(3), sum(2) => SUM(2), sum(1) => SUM(1), sum(0) 
                           => SUM(0));
   SBi_1 : SUM_BLOCK_K4_7 port map( a(3) => A(7), a(2) => A(6), a(1) => A(5), 
                           a(0) => A(4), b(3) => B(7), b(2) => B(6), b(1) => 
                           B(5), b(0) => B(4), C_gen => carries(1), sum(3) => 
                           SUM(7), sum(2) => SUM(6), sum(1) => SUM(5), sum(0) 
                           => SUM(4));
   SBi_2 : SUM_BLOCK_K4_6 port map( a(3) => A(11), a(2) => A(10), a(1) => A(9),
                           a(0) => A(8), b(3) => B(11), b(2) => B(10), b(1) => 
                           B(9), b(0) => B(8), C_gen => carries(2), sum(3) => 
                           SUM(11), sum(2) => SUM(10), sum(1) => SUM(9), sum(0)
                           => SUM(8));
   SBi_3 : SUM_BLOCK_K4_5 port map( a(3) => A(15), a(2) => A(14), a(1) => A(13)
                           , a(0) => A(12), b(3) => B(15), b(2) => B(14), b(1) 
                           => B(13), b(0) => B(12), C_gen => carries(3), sum(3)
                           => SUM(15), sum(2) => SUM(14), sum(1) => SUM(13), 
                           sum(0) => SUM(12));
   SBi_4 : SUM_BLOCK_K4_4 port map( a(3) => A(19), a(2) => A(18), a(1) => A(17)
                           , a(0) => A(16), b(3) => B(19), b(2) => B(18), b(1) 
                           => B(17), b(0) => B(16), C_gen => carries(4), sum(3)
                           => SUM(19), sum(2) => SUM(18), sum(1) => SUM(17), 
                           sum(0) => SUM(16));
   SBi_5 : SUM_BLOCK_K4_3 port map( a(3) => A(23), a(2) => A(22), a(1) => A(21)
                           , a(0) => A(20), b(3) => B(23), b(2) => B(22), b(1) 
                           => B(21), b(0) => B(20), C_gen => carries(5), sum(3)
                           => SUM(23), sum(2) => SUM(22), sum(1) => SUM(21), 
                           sum(0) => SUM(20));
   SBi_6 : SUM_BLOCK_K4_2 port map( a(3) => A(27), a(2) => A(26), a(1) => A(25)
                           , a(0) => A(24), b(3) => B(27), b(2) => B(26), b(1) 
                           => B(25), b(0) => B(24), C_gen => carries(6), sum(3)
                           => SUM(27), sum(2) => SUM(26), sum(1) => SUM(25), 
                           sum(0) => SUM(24));
   SBi_7 : SUM_BLOCK_K4_1 port map( a(3) => A(31), a(2) => A(30), a(1) => A(29)
                           , a(0) => A(28), b(3) => B(31), b(2) => B(30), b(1) 
                           => B(29), b(0) => B(28), C_gen => carries(7), sum(3)
                           => SUM(31), sum(2) => SUM(30), sum(1) => SUM(29), 
                           sum(0) => SUM(28));

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity CARRY_GENERATOR_NBIT32_NBLOCK4 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co : 
         out std_logic_vector (8 downto 0));

end CARRY_GENERATOR_NBIT32_NBLOCK4;

architecture SYN_Structural of CARRY_GENERATOR_NBIT32_NBLOCK4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component G_BLOCK_1
      port( PIK, GIK, GK1J : in std_logic;  GIJ : out std_logic);
   end component;
   
   component G_BLOCK_2
      port( PIK, GIK, GK1J : in std_logic;  GIJ : out std_logic);
   end component;
   
   component G_BLOCK_3
      port( PIK, GIK, GK1J : in std_logic;  GIJ : out std_logic);
   end component;
   
   component G_BLOCK_4
      port( PIK, GIK, GK1J : in std_logic;  GIJ : out std_logic);
   end component;
   
   component PG_BLOCK_1
      port( PIK, GIK, PK1J, GK1J : in std_logic;  GIJ, PIJ : out std_logic);
   end component;
   
   component PG_BLOCK_2
      port( PIK, GIK, PK1J, GK1J : in std_logic;  GIJ, PIJ : out std_logic);
   end component;
   
   component G_BLOCK_5
      port( PIK, GIK, GK1J : in std_logic;  GIJ : out std_logic);
   end component;
   
   component G_BLOCK_6
      port( PIK, GIK, GK1J : in std_logic;  GIJ : out std_logic);
   end component;
   
   component PG_BLOCK_3
      port( PIK, GIK, PK1J, GK1J : in std_logic;  GIJ, PIJ : out std_logic);
   end component;
   
   component PG_BLOCK_4
      port( PIK, GIK, PK1J, GK1J : in std_logic;  GIJ, PIJ : out std_logic);
   end component;
   
   component PG_BLOCK_5
      port( PIK, GIK, PK1J, GK1J : in std_logic;  GIJ, PIJ : out std_logic);
   end component;
   
   component G_BLOCK_7
      port( PIK, GIK, GK1J : in std_logic;  GIJ : out std_logic);
   end component;
   
   component PG_BLOCK_6
      port( PIK, GIK, PK1J, GK1J : in std_logic;  GIJ, PIJ : out std_logic);
   end component;
   
   component PG_BLOCK_7
      port( PIK, GIK, PK1J, GK1J : in std_logic;  GIJ, PIJ : out std_logic);
   end component;
   
   component PG_BLOCK_8
      port( PIK, GIK, PK1J, GK1J : in std_logic;  GIJ, PIJ : out std_logic);
   end component;
   
   component PG_BLOCK_9
      port( PIK, GIK, PK1J, GK1J : in std_logic;  GIJ, PIJ : out std_logic);
   end component;
   
   component PG_BLOCK_10
      port( PIK, GIK, PK1J, GK1J : in std_logic;  GIJ, PIJ : out std_logic);
   end component;
   
   component PG_BLOCK_11
      port( PIK, GIK, PK1J, GK1J : in std_logic;  GIJ, PIJ : out std_logic);
   end component;
   
   component PG_BLOCK_12
      port( PIK, GIK, PK1J, GK1J : in std_logic;  GIJ, PIJ : out std_logic);
   end component;
   
   component G_BLOCK_8
      port( PIK, GIK, GK1J : in std_logic;  GIJ : out std_logic);
   end component;
   
   component PG_BLOCK_13
      port( PIK, GIK, PK1J, GK1J : in std_logic;  GIJ, PIJ : out std_logic);
   end component;
   
   component PG_BLOCK_14
      port( PIK, GIK, PK1J, GK1J : in std_logic;  GIJ, PIJ : out std_logic);
   end component;
   
   component PG_BLOCK_15
      port( PIK, GIK, PK1J, GK1J : in std_logic;  GIJ, PIJ : out std_logic);
   end component;
   
   component PG_BLOCK_16
      port( PIK, GIK, PK1J, GK1J : in std_logic;  GIJ, PIJ : out std_logic);
   end component;
   
   component PG_BLOCK_17
      port( PIK, GIK, PK1J, GK1J : in std_logic;  GIJ, PIJ : out std_logic);
   end component;
   
   component PG_BLOCK_18
      port( PIK, GIK, PK1J, GK1J : in std_logic;  GIJ, PIJ : out std_logic);
   end component;
   
   component PG_BLOCK_19
      port( PIK, GIK, PK1J, GK1J : in std_logic;  GIJ, PIJ : out std_logic);
   end component;
   
   component PG_BLOCK_20
      port( PIK, GIK, PK1J, GK1J : in std_logic;  GIJ, PIJ : out std_logic);
   end component;
   
   component PG_BLOCK_21
      port( PIK, GIK, PK1J, GK1J : in std_logic;  GIJ, PIJ : out std_logic);
   end component;
   
   component PG_BLOCK_22
      port( PIK, GIK, PK1J, GK1J : in std_logic;  GIJ, PIJ : out std_logic);
   end component;
   
   component PG_BLOCK_23
      port( PIK, GIK, PK1J, GK1J : in std_logic;  GIJ, PIJ : out std_logic);
   end component;
   
   component PG_BLOCK_24
      port( PIK, GIK, PK1J, GK1J : in std_logic;  GIJ, PIJ : out std_logic);
   end component;
   
   component PG_BLOCK_25
      port( PIK, GIK, PK1J, GK1J : in std_logic;  GIJ, PIJ : out std_logic);
   end component;
   
   component PG_BLOCK_26
      port( PIK, GIK, PK1J, GK1J : in std_logic;  GIJ, PIJ : out std_logic);
   end component;
   
   component PG_BLOCK_0
      port( PIK, GIK, PK1J, GK1J : in std_logic;  GIJ, PIJ : out std_logic);
   end component;
   
   component G_BLOCK_0
      port( PIK, GIK, GK1J : in std_logic;  GIJ : out std_logic);
   end component;
   
   component PG_NET_1
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_NET_2
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_NET_3
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_NET_4
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_NET_5
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_NET_6
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_NET_7
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_NET_8
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_NET_9
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_NET_10
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_NET_11
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_NET_12
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_NET_13
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_NET_14
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_NET_15
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_NET_16
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_NET_17
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_NET_18
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_NET_19
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_NET_20
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_NET_21
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_NET_22
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_NET_23
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_NET_24
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_NET_25
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_NET_26
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_NET_27
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_NET_28
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_NET_29
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_NET_30
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_NET_31
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_NET_0
      port( A, B : in std_logic;  P, G : out std_logic);
   end component;
   
   signal Co_8_port, Co_7_port, Co_6_port, Co_5_port, n8, Co_3_port, n9, n10, 
      PGNET_G_4_31_port, PGNET_G_4_27_port, PGNET_G_3_31_port, 
      PGNET_G_3_23_port, PGNET_G_3_15_port, PGNET_G_3_11_port, 
      PGNET_G_2_31_port, PGNET_G_2_27_port, PGNET_G_2_23_port, 
      PGNET_G_2_19_port, PGNET_G_2_15_port, PGNET_G_2_7_port, PGNET_G_1_31_port
      , PGNET_G_1_29_port, PGNET_G_1_27_port, PGNET_G_1_25_port, 
      PGNET_G_1_23_port, PGNET_G_1_21_port, PGNET_G_1_19_port, 
      PGNET_G_1_17_port, PGNET_G_1_15_port, PGNET_G_1_13_port, 
      PGNET_G_1_11_port, PGNET_G_1_9_port, PGNET_G_1_7_port, PGNET_G_1_5_port, 
      PGNET_G_1_3_port, PGNET_G_0_31_port, PGNET_G_0_30_port, PGNET_G_0_29_port
      , PGNET_G_0_28_port, PGNET_G_0_27_port, PGNET_G_0_26_port, 
      PGNET_G_0_25_port, PGNET_G_0_24_port, PGNET_G_0_23_port, 
      PGNET_G_0_22_port, PGNET_G_0_21_port, PGNET_G_0_20_port, 
      PGNET_G_0_19_port, PGNET_G_0_18_port, PGNET_G_0_17_port, 
      PGNET_G_0_16_port, PGNET_G_0_15_port, PGNET_G_0_14_port, 
      PGNET_G_0_13_port, PGNET_G_0_12_port, PGNET_G_0_11_port, 
      PGNET_G_0_10_port, PGNET_G_0_9_port, PGNET_G_0_8_port, PGNET_G_0_7_port, 
      PGNET_G_0_6_port, PGNET_G_0_5_port, PGNET_G_0_4_port, PGNET_G_0_3_port, 
      PGNET_G_0_2_port, PGNET_G_0_1_port, PGNET_G_0_0_port, PGNET_P_4_31_port, 
      PGNET_P_4_27_port, PGNET_P_3_31_port, PGNET_P_3_23_port, 
      PGNET_P_3_15_port, PGNET_P_3_11_port, PGNET_P_2_31_port, 
      PGNET_P_2_27_port, PGNET_P_2_23_port, PGNET_P_2_19_port, 
      PGNET_P_2_15_port, PGNET_P_2_7_port, PGNET_P_1_31_port, PGNET_P_1_29_port
      , PGNET_P_1_27_port, PGNET_P_1_25_port, PGNET_P_1_23_port, 
      PGNET_P_1_21_port, PGNET_P_1_19_port, PGNET_P_1_17_port, 
      PGNET_P_1_15_port, PGNET_P_1_13_port, PGNET_P_1_11_port, PGNET_P_1_9_port
      , PGNET_P_1_7_port, PGNET_P_1_5_port, PGNET_P_1_3_port, PGNET_P_0_31_port
      , PGNET_P_0_30_port, PGNET_P_0_29_port, PGNET_P_0_28_port, 
      PGNET_P_0_27_port, PGNET_P_0_26_port, PGNET_P_0_25_port, 
      PGNET_P_0_24_port, PGNET_P_0_23_port, PGNET_P_0_22_port, 
      PGNET_P_0_21_port, PGNET_P_0_20_port, PGNET_P_0_19_port, 
      PGNET_P_0_18_port, PGNET_P_0_17_port, PGNET_P_0_16_port, 
      PGNET_P_0_15_port, PGNET_P_0_14_port, PGNET_P_0_13_port, 
      PGNET_P_0_12_port, PGNET_P_0_11_port, PGNET_P_0_10_port, PGNET_P_0_9_port
      , PGNET_P_0_8_port, PGNET_P_0_7_port, PGNET_P_0_6_port, PGNET_P_0_5_port,
      PGNET_P_0_4_port, PGNET_P_0_3_port, PGNET_P_0_2_port, PGNET_P_0_1_port, 
      carries_1_port, n11, n12, Co_4_port, n14, Co_1_port, n16, Co_2_port, 
      n_1016 : std_logic;

begin
   Co <= ( Co_8_port, Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, 
      Co_2_port, Co_1_port, Cin );
   
   pgport_0 : PG_NET_0 port map( A => A(0), B => B(0), P => n_1016, G => 
                           PGNET_G_0_0_port);
   pgport_1 : PG_NET_31 port map( A => A(1), B => B(1), P => PGNET_P_0_1_port, 
                           G => PGNET_G_0_1_port);
   pgport_2 : PG_NET_30 port map( A => A(2), B => B(2), P => PGNET_P_0_2_port, 
                           G => PGNET_G_0_2_port);
   pgport_3 : PG_NET_29 port map( A => A(3), B => B(3), P => PGNET_P_0_3_port, 
                           G => PGNET_G_0_3_port);
   pgport_4 : PG_NET_28 port map( A => A(4), B => B(4), P => PGNET_P_0_4_port, 
                           G => PGNET_G_0_4_port);
   pgport_5 : PG_NET_27 port map( A => A(5), B => B(5), P => PGNET_P_0_5_port, 
                           G => PGNET_G_0_5_port);
   pgport_6 : PG_NET_26 port map( A => A(6), B => B(6), P => PGNET_P_0_6_port, 
                           G => PGNET_G_0_6_port);
   pgport_7 : PG_NET_25 port map( A => A(7), B => B(7), P => PGNET_P_0_7_port, 
                           G => PGNET_G_0_7_port);
   pgport_8 : PG_NET_24 port map( A => A(8), B => B(8), P => PGNET_P_0_8_port, 
                           G => PGNET_G_0_8_port);
   pgport_9 : PG_NET_23 port map( A => A(9), B => B(9), P => PGNET_P_0_9_port, 
                           G => PGNET_G_0_9_port);
   pgport_10 : PG_NET_22 port map( A => A(10), B => B(10), P => 
                           PGNET_P_0_10_port, G => PGNET_G_0_10_port);
   pgport_11 : PG_NET_21 port map( A => A(11), B => B(11), P => 
                           PGNET_P_0_11_port, G => PGNET_G_0_11_port);
   pgport_12 : PG_NET_20 port map( A => A(12), B => B(12), P => 
                           PGNET_P_0_12_port, G => PGNET_G_0_12_port);
   pgport_13 : PG_NET_19 port map( A => A(13), B => B(13), P => 
                           PGNET_P_0_13_port, G => PGNET_G_0_13_port);
   pgport_14 : PG_NET_18 port map( A => A(14), B => B(14), P => 
                           PGNET_P_0_14_port, G => PGNET_G_0_14_port);
   pgport_15 : PG_NET_17 port map( A => A(15), B => B(15), P => 
                           PGNET_P_0_15_port, G => PGNET_G_0_15_port);
   pgport_16 : PG_NET_16 port map( A => A(16), B => B(16), P => 
                           PGNET_P_0_16_port, G => PGNET_G_0_16_port);
   pgport_17 : PG_NET_15 port map( A => A(17), B => B(17), P => 
                           PGNET_P_0_17_port, G => PGNET_G_0_17_port);
   pgport_18 : PG_NET_14 port map( A => A(18), B => B(18), P => 
                           PGNET_P_0_18_port, G => PGNET_G_0_18_port);
   pgport_19 : PG_NET_13 port map( A => A(19), B => B(19), P => 
                           PGNET_P_0_19_port, G => PGNET_G_0_19_port);
   pgport_20 : PG_NET_12 port map( A => A(20), B => B(20), P => 
                           PGNET_P_0_20_port, G => PGNET_G_0_20_port);
   pgport_21 : PG_NET_11 port map( A => A(21), B => B(21), P => 
                           PGNET_P_0_21_port, G => PGNET_G_0_21_port);
   pgport_22 : PG_NET_10 port map( A => A(22), B => B(22), P => 
                           PGNET_P_0_22_port, G => PGNET_G_0_22_port);
   pgport_23 : PG_NET_9 port map( A => A(23), B => B(23), P => 
                           PGNET_P_0_23_port, G => PGNET_G_0_23_port);
   pgport_24 : PG_NET_8 port map( A => A(24), B => B(24), P => 
                           PGNET_P_0_24_port, G => PGNET_G_0_24_port);
   pgport_25 : PG_NET_7 port map( A => A(25), B => B(25), P => 
                           PGNET_P_0_25_port, G => PGNET_G_0_25_port);
   pgport_26 : PG_NET_6 port map( A => A(26), B => B(26), P => 
                           PGNET_P_0_26_port, G => PGNET_G_0_26_port);
   pgport_27 : PG_NET_5 port map( A => A(27), B => B(27), P => 
                           PGNET_P_0_27_port, G => PGNET_G_0_27_port);
   pgport_28 : PG_NET_4 port map( A => A(28), B => B(28), P => 
                           PGNET_P_0_28_port, G => PGNET_G_0_28_port);
   pgport_29 : PG_NET_3 port map( A => A(29), B => B(29), P => 
                           PGNET_P_0_29_port, G => PGNET_G_0_29_port);
   pgport_30 : PG_NET_2 port map( A => A(30), B => B(30), P => 
                           PGNET_P_0_30_port, G => PGNET_G_0_30_port);
   pgport_31 : PG_NET_1 port map( A => A(31), B => B(31), P => 
                           PGNET_P_0_31_port, G => PGNET_G_0_31_port);
   gi_1_1 : G_BLOCK_0 port map( PIK => PGNET_P_0_1_port, GIK => 
                           PGNET_G_0_1_port, GK1J => PGNET_G_0_0_port, GIJ => 
                           carries_1_port);
   pgi_1_3 : PG_BLOCK_0 port map( PIK => PGNET_P_0_3_port, GIK => 
                           PGNET_G_0_3_port, PK1J => PGNET_P_0_2_port, GK1J => 
                           PGNET_G_0_2_port, GIJ => PGNET_G_1_3_port, PIJ => 
                           PGNET_P_1_3_port);
   pgi_1_5 : PG_BLOCK_26 port map( PIK => PGNET_P_0_5_port, GIK => 
                           PGNET_G_0_5_port, PK1J => PGNET_P_0_4_port, GK1J => 
                           PGNET_G_0_4_port, GIJ => PGNET_G_1_5_port, PIJ => 
                           PGNET_P_1_5_port);
   pgi_1_7 : PG_BLOCK_25 port map( PIK => PGNET_P_0_7_port, GIK => 
                           PGNET_G_0_7_port, PK1J => PGNET_P_0_6_port, GK1J => 
                           PGNET_G_0_6_port, GIJ => PGNET_G_1_7_port, PIJ => 
                           PGNET_P_1_7_port);
   pgi_1_9 : PG_BLOCK_24 port map( PIK => PGNET_P_0_9_port, GIK => 
                           PGNET_G_0_9_port, PK1J => PGNET_P_0_8_port, GK1J => 
                           PGNET_G_0_8_port, GIJ => PGNET_G_1_9_port, PIJ => 
                           PGNET_P_1_9_port);
   pgi_1_11 : PG_BLOCK_23 port map( PIK => PGNET_P_0_11_port, GIK => 
                           PGNET_G_0_11_port, PK1J => PGNET_P_0_10_port, GK1J 
                           => PGNET_G_0_10_port, GIJ => PGNET_G_1_11_port, PIJ 
                           => PGNET_P_1_11_port);
   pgi_1_13 : PG_BLOCK_22 port map( PIK => PGNET_P_0_13_port, GIK => 
                           PGNET_G_0_13_port, PK1J => PGNET_P_0_12_port, GK1J 
                           => PGNET_G_0_12_port, GIJ => PGNET_G_1_13_port, PIJ 
                           => PGNET_P_1_13_port);
   pgi_1_15 : PG_BLOCK_21 port map( PIK => PGNET_P_0_15_port, GIK => 
                           PGNET_G_0_15_port, PK1J => PGNET_P_0_14_port, GK1J 
                           => PGNET_G_0_14_port, GIJ => PGNET_G_1_15_port, PIJ 
                           => PGNET_P_1_15_port);
   pgi_1_17 : PG_BLOCK_20 port map( PIK => PGNET_P_0_17_port, GIK => 
                           PGNET_G_0_17_port, PK1J => PGNET_P_0_16_port, GK1J 
                           => PGNET_G_0_16_port, GIJ => PGNET_G_1_17_port, PIJ 
                           => PGNET_P_1_17_port);
   pgi_1_19 : PG_BLOCK_19 port map( PIK => PGNET_P_0_19_port, GIK => 
                           PGNET_G_0_19_port, PK1J => PGNET_P_0_18_port, GK1J 
                           => PGNET_G_0_18_port, GIJ => PGNET_G_1_19_port, PIJ 
                           => PGNET_P_1_19_port);
   pgi_1_21 : PG_BLOCK_18 port map( PIK => PGNET_P_0_21_port, GIK => 
                           PGNET_G_0_21_port, PK1J => PGNET_P_0_20_port, GK1J 
                           => PGNET_G_0_20_port, GIJ => PGNET_G_1_21_port, PIJ 
                           => PGNET_P_1_21_port);
   pgi_1_23 : PG_BLOCK_17 port map( PIK => PGNET_P_0_23_port, GIK => 
                           PGNET_G_0_23_port, PK1J => PGNET_P_0_22_port, GK1J 
                           => PGNET_G_0_22_port, GIJ => PGNET_G_1_23_port, PIJ 
                           => PGNET_P_1_23_port);
   pgi_1_25 : PG_BLOCK_16 port map( PIK => PGNET_P_0_25_port, GIK => 
                           PGNET_G_0_25_port, PK1J => PGNET_P_0_24_port, GK1J 
                           => PGNET_G_0_24_port, GIJ => PGNET_G_1_25_port, PIJ 
                           => PGNET_P_1_25_port);
   pgi_1_27 : PG_BLOCK_15 port map( PIK => PGNET_P_0_27_port, GIK => 
                           PGNET_G_0_27_port, PK1J => PGNET_P_0_26_port, GK1J 
                           => PGNET_G_0_26_port, GIJ => PGNET_G_1_27_port, PIJ 
                           => PGNET_P_1_27_port);
   pgi_1_29 : PG_BLOCK_14 port map( PIK => PGNET_P_0_29_port, GIK => 
                           PGNET_G_0_29_port, PK1J => PGNET_P_0_28_port, GK1J 
                           => PGNET_G_0_28_port, GIJ => PGNET_G_1_29_port, PIJ 
                           => PGNET_P_1_29_port);
   pgi_1_31 : PG_BLOCK_13 port map( PIK => PGNET_P_0_31_port, GIK => 
                           PGNET_G_0_31_port, PK1J => PGNET_P_0_30_port, GK1J 
                           => PGNET_G_0_30_port, GIJ => PGNET_G_1_31_port, PIJ 
                           => PGNET_P_1_31_port);
   gi_2_3 : G_BLOCK_8 port map( PIK => PGNET_P_1_3_port, GIK => 
                           PGNET_G_1_3_port, GK1J => carries_1_port, GIJ => n10
                           );
   pgi_2_7 : PG_BLOCK_12 port map( PIK => PGNET_P_1_7_port, GIK => 
                           PGNET_G_1_7_port, PK1J => PGNET_P_1_5_port, GK1J => 
                           PGNET_G_1_5_port, GIJ => PGNET_G_2_7_port, PIJ => 
                           PGNET_P_2_7_port);
   pgi_2_11 : PG_BLOCK_11 port map( PIK => PGNET_P_1_11_port, GIK => 
                           PGNET_G_1_11_port, PK1J => PGNET_P_1_9_port, GK1J =>
                           PGNET_G_1_9_port, GIJ => PGNET_G_3_11_port, PIJ => 
                           PGNET_P_3_11_port);
   pgi_2_15 : PG_BLOCK_10 port map( PIK => PGNET_P_1_15_port, GIK => 
                           PGNET_G_1_15_port, PK1J => PGNET_P_1_13_port, GK1J 
                           => PGNET_G_1_13_port, GIJ => PGNET_G_2_15_port, PIJ 
                           => PGNET_P_2_15_port);
   pgi_2_19 : PG_BLOCK_9 port map( PIK => PGNET_P_1_19_port, GIK => 
                           PGNET_G_1_19_port, PK1J => PGNET_P_1_17_port, GK1J 
                           => PGNET_G_1_17_port, GIJ => PGNET_G_2_19_port, PIJ 
                           => PGNET_P_2_19_port);
   pgi_2_23 : PG_BLOCK_8 port map( PIK => PGNET_P_1_23_port, GIK => 
                           PGNET_G_1_23_port, PK1J => PGNET_P_1_21_port, GK1J 
                           => PGNET_G_1_21_port, GIJ => PGNET_G_2_23_port, PIJ 
                           => PGNET_P_2_23_port);
   pgi_2_27 : PG_BLOCK_7 port map( PIK => PGNET_P_1_27_port, GIK => 
                           PGNET_G_1_27_port, PK1J => PGNET_P_1_25_port, GK1J 
                           => PGNET_G_1_25_port, GIJ => PGNET_G_2_27_port, PIJ 
                           => PGNET_P_2_27_port);
   pgi_2_31 : PG_BLOCK_6 port map( PIK => PGNET_P_1_31_port, GIK => 
                           PGNET_G_1_31_port, PK1J => PGNET_P_1_29_port, GK1J 
                           => PGNET_G_1_29_port, GIJ => PGNET_G_2_31_port, PIJ 
                           => PGNET_P_2_31_port);
   gi_3_7 : G_BLOCK_7 port map( PIK => PGNET_P_2_7_port, GIK => 
                           PGNET_G_2_7_port, GK1J => n10, GIJ => n9);
   pgi_3_15 : PG_BLOCK_5 port map( PIK => PGNET_P_2_15_port, GIK => 
                           PGNET_G_2_15_port, PK1J => PGNET_P_3_11_port, GK1J 
                           => PGNET_G_3_11_port, GIJ => PGNET_G_3_15_port, PIJ 
                           => PGNET_P_3_15_port);
   pgi_3_23 : PG_BLOCK_4 port map( PIK => PGNET_P_2_23_port, GIK => 
                           PGNET_G_2_23_port, PK1J => PGNET_P_2_19_port, GK1J 
                           => PGNET_G_2_19_port, GIJ => PGNET_G_3_23_port, PIJ 
                           => PGNET_P_3_23_port);
   pgi_3_31 : PG_BLOCK_3 port map( PIK => PGNET_P_2_31_port, GIK => 
                           PGNET_G_2_31_port, PK1J => PGNET_P_2_27_port, GK1J 
                           => PGNET_G_2_27_port, GIJ => PGNET_G_3_31_port, PIJ 
                           => PGNET_P_3_31_port);
   gi_4_11 : G_BLOCK_6 port map( PIK => PGNET_P_3_11_port, GIK => 
                           PGNET_G_3_11_port, GK1J => n12, GIJ => Co_3_port);
   gi_4_15 : G_BLOCK_5 port map( PIK => PGNET_P_3_15_port, GIK => 
                           PGNET_G_3_15_port, GK1J => n9, GIJ => n8);
   pgi_4_27 : PG_BLOCK_2 port map( PIK => PGNET_P_2_27_port, GIK => 
                           PGNET_G_2_27_port, PK1J => PGNET_P_3_23_port, GK1J 
                           => PGNET_G_3_23_port, GIJ => PGNET_G_4_27_port, PIJ 
                           => PGNET_P_4_27_port);
   pgi_4_31 : PG_BLOCK_1 port map( PIK => PGNET_P_3_31_port, GIK => 
                           PGNET_G_3_31_port, PK1J => PGNET_P_3_23_port, GK1J 
                           => n11, GIJ => PGNET_G_4_31_port, PIJ => 
                           PGNET_P_4_31_port);
   gi_5_19 : G_BLOCK_4 port map( PIK => PGNET_P_2_19_port, GIK => 
                           PGNET_G_2_19_port, GK1J => n8, GIJ => Co_5_port);
   gi_5_23 : G_BLOCK_3 port map( PIK => PGNET_P_3_23_port, GIK => n11, GK1J => 
                           n8, GIJ => Co_6_port);
   gi_5_27 : G_BLOCK_2 port map( PIK => PGNET_P_4_27_port, GIK => 
                           PGNET_G_4_27_port, GK1J => n8, GIJ => Co_7_port);
   gi_5_31 : G_BLOCK_1 port map( PIK => PGNET_P_4_31_port, GIK => 
                           PGNET_G_4_31_port, GK1J => Co_4_port, GIJ => 
                           Co_8_port);
   U1 : CLKBUF_X1 port map( A => PGNET_G_3_23_port, Z => n11);
   U2 : INV_X1 port map( A => n16, ZN => n12);
   U3 : BUF_X2 port map( A => n14, Z => Co_4_port);
   U4 : CLKBUF_X1 port map( A => n8, Z => n14);
   U5 : CLKBUF_X1 port map( A => n10, Z => Co_1_port);
   U6 : INV_X1 port map( A => n9, ZN => n16);
   U7 : INV_X1 port map( A => n16, ZN => Co_2_port);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4Adder.all;

entity P4Adder is

   port( A, B : in std_logic_vector (31 downto 0);  CIN : in std_logic;  Cout :
         out std_logic;  SUM : out std_logic_vector (31 downto 0));

end P4Adder;

architecture SYN_Structural of P4Adder is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component SUM_GENERATOR_N32_K4
      port( carries : in std_logic_vector (7 downto 0);  A, B : in 
            std_logic_vector (31 downto 0);  SUM : out std_logic_vector (31 
            downto 0));
   end component;
   
   component CARRY_GENERATOR_NBIT32_NBLOCK4
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co 
            : out std_logic_vector (8 downto 0));
   end component;
   
   signal carries_s_7_port, carries_s_6_port, carries_s_5_port, 
      carries_s_4_port, carries_s_3_port, carries_s_2_port, carries_s_1_port, 
      carries_s_0_port, n1, n2, n3, n4 : std_logic;

begin
   
   CG : CARRY_GENERATOR_NBIT32_NBLOCK4 port map( A(31) => A(31), A(30) => A(30)
                           , A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Cin => CIN, Co(8) => Cout, Co(7)
                           => carries_s_7_port, Co(6) => carries_s_6_port, 
                           Co(5) => carries_s_5_port, Co(4) => carries_s_4_port
                           , Co(3) => carries_s_3_port, Co(2) => 
                           carries_s_2_port, Co(1) => carries_s_1_port, Co(0) 
                           => carries_s_0_port);
   SG : SUM_GENERATOR_N32_K4 port map( carries(7) => carries_s_7_port, 
                           carries(6) => carries_s_6_port, carries(5) => 
                           carries_s_5_port, carries(4) => carries_s_4_port, 
                           carries(3) => carries_s_3_port, carries(2) => 
                           carries_s_2_port, carries(1) => carries_s_1_port, 
                           carries(0) => carries_s_0_port, A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => n2, A(14) => A(14), A(13) => A(13), A(12) 
                           => A(12), A(11) => A(11), A(10) => A(10), A(9) => 
                           A(9), A(8) => A(8), A(7) => n4, A(6) => A(6), A(5) 
                           => A(5), A(4) => A(4), A(3) => n3, A(2) => A(2), 
                           A(1) => A(1), A(0) => A(0), B(31) => B(31), B(30) =>
                           B(30), B(29) => B(29), B(28) => B(28), B(27) => 
                           B(27), B(26) => B(26), B(25) => B(25), B(24) => 
                           B(24), B(23) => B(23), B(22) => B(22), B(21) => 
                           B(21), B(20) => B(20), B(19) => B(19), B(18) => 
                           B(18), B(17) => B(17), B(16) => B(16), B(15) => n1, 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), SUM(31) => SUM(31), SUM(30) => 
                           SUM(30), SUM(29) => SUM(29), SUM(28) => SUM(28), 
                           SUM(27) => SUM(27), SUM(26) => SUM(26), SUM(25) => 
                           SUM(25), SUM(24) => SUM(24), SUM(23) => SUM(23), 
                           SUM(22) => SUM(22), SUM(21) => SUM(21), SUM(20) => 
                           SUM(20), SUM(19) => SUM(19), SUM(18) => SUM(18), 
                           SUM(17) => SUM(17), SUM(16) => SUM(16), SUM(15) => 
                           SUM(15), SUM(14) => SUM(14), SUM(13) => SUM(13), 
                           SUM(12) => SUM(12), SUM(11) => SUM(11), SUM(10) => 
                           SUM(10), SUM(9) => SUM(9), SUM(8) => SUM(8), SUM(7) 
                           => SUM(7), SUM(6) => SUM(6), SUM(5) => SUM(5), 
                           SUM(4) => SUM(4), SUM(3) => SUM(3), SUM(2) => SUM(2)
                           , SUM(1) => SUM(1), SUM(0) => SUM(0));
   U1 : BUF_X1 port map( A => B(15), Z => n1);
   U2 : BUF_X1 port map( A => A(15), Z => n2);
   U3 : BUF_X1 port map( A => A(3), Z => n3);
   U4 : BUF_X1 port map( A => A(7), Z => n4);

end SYN_Structural;
